module Swapper(
  input  [7:0] io_a0,
  input  [7:0] io_a1,
  output [7:0] io_z0,
  output [7:0] io_z1
);
  wire  _T; // @[bitonic_sort.scala 62:89]
  assign _T = io_a1 < io_a0; // @[bitonic_sort.scala 62:89]
  assign io_z0 = _T ? io_a1 : io_a0; // @[bitonic_sort.scala 15:11 bitonic_sort.scala 18:11]
  assign io_z1 = _T ? io_a0 : io_a1; // @[bitonic_sort.scala 16:11 bitonic_sort.scala 19:11]
endmodule
module BitonicSorterModule(
  input        clock,
  input        reset,
  input  [7:0] io_a_0,
  input  [7:0] io_a_1,
  input  [7:0] io_a_2,
  input  [7:0] io_a_3,
  input  [7:0] io_a_4,
  input  [7:0] io_a_5,
  input  [7:0] io_a_6,
  input  [7:0] io_a_7,
  input  [7:0] io_a_8,
  input  [7:0] io_a_9,
  input  [7:0] io_a_10,
  input  [7:0] io_a_11,
  input  [7:0] io_a_12,
  input  [7:0] io_a_13,
  input  [7:0] io_a_14,
  input  [7:0] io_a_15,
  input  [7:0] io_a_16,
  input  [7:0] io_a_17,
  input  [7:0] io_a_18,
  input  [7:0] io_a_19,
  input  [7:0] io_a_20,
  input  [7:0] io_a_21,
  input  [7:0] io_a_22,
  input  [7:0] io_a_23,
  input  [7:0] io_a_24,
  input  [7:0] io_a_25,
  input  [7:0] io_a_26,
  input  [7:0] io_a_27,
  input  [7:0] io_a_28,
  input  [7:0] io_a_29,
  input  [7:0] io_a_30,
  input  [7:0] io_a_31,
  input  [7:0] io_a_32,
  input  [7:0] io_a_33,
  input  [7:0] io_a_34,
  input  [7:0] io_a_35,
  input  [7:0] io_a_36,
  input  [7:0] io_a_37,
  input  [7:0] io_a_38,
  input  [7:0] io_a_39,
  input  [7:0] io_a_40,
  input  [7:0] io_a_41,
  input  [7:0] io_a_42,
  input  [7:0] io_a_43,
  input  [7:0] io_a_44,
  input  [7:0] io_a_45,
  input  [7:0] io_a_46,
  input  [7:0] io_a_47,
  input  [7:0] io_a_48,
  input  [7:0] io_a_49,
  input  [7:0] io_a_50,
  input  [7:0] io_a_51,
  input  [7:0] io_a_52,
  input  [7:0] io_a_53,
  input  [7:0] io_a_54,
  input  [7:0] io_a_55,
  input  [7:0] io_a_56,
  input  [7:0] io_a_57,
  input  [7:0] io_a_58,
  input  [7:0] io_a_59,
  input  [7:0] io_a_60,
  input  [7:0] io_a_61,
  input  [7:0] io_a_62,
  input  [7:0] io_a_63,
  output [7:0] io_z_0,
  output [7:0] io_z_1,
  output [7:0] io_z_2,
  output [7:0] io_z_3,
  output [7:0] io_z_4,
  output [7:0] io_z_5,
  output [7:0] io_z_6,
  output [7:0] io_z_7,
  output [7:0] io_z_8,
  output [7:0] io_z_9,
  output [7:0] io_z_10,
  output [7:0] io_z_11,
  output [7:0] io_z_12,
  output [7:0] io_z_13,
  output [7:0] io_z_14,
  output [7:0] io_z_15,
  output [7:0] io_z_16,
  output [7:0] io_z_17,
  output [7:0] io_z_18,
  output [7:0] io_z_19,
  output [7:0] io_z_20,
  output [7:0] io_z_21,
  output [7:0] io_z_22,
  output [7:0] io_z_23,
  output [7:0] io_z_24,
  output [7:0] io_z_25,
  output [7:0] io_z_26,
  output [7:0] io_z_27,
  output [7:0] io_z_28,
  output [7:0] io_z_29,
  output [7:0] io_z_30,
  output [7:0] io_z_31,
  output [7:0] io_z_32,
  output [7:0] io_z_33,
  output [7:0] io_z_34,
  output [7:0] io_z_35,
  output [7:0] io_z_36,
  output [7:0] io_z_37,
  output [7:0] io_z_38,
  output [7:0] io_z_39,
  output [7:0] io_z_40,
  output [7:0] io_z_41,
  output [7:0] io_z_42,
  output [7:0] io_z_43,
  output [7:0] io_z_44,
  output [7:0] io_z_45,
  output [7:0] io_z_46,
  output [7:0] io_z_47,
  output [7:0] io_z_48,
  output [7:0] io_z_49,
  output [7:0] io_z_50,
  output [7:0] io_z_51,
  output [7:0] io_z_52,
  output [7:0] io_z_53,
  output [7:0] io_z_54,
  output [7:0] io_z_55,
  output [7:0] io_z_56,
  output [7:0] io_z_57,
  output [7:0] io_z_58,
  output [7:0] io_z_59,
  output [7:0] io_z_60,
  output [7:0] io_z_61,
  output [7:0] io_z_62,
  output [7:0] io_z_63
);
  wire [7:0] Swapper_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_1_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_1_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_1_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_1_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_2_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_2_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_2_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_2_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_3_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_3_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_3_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_3_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_4_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_4_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_4_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_4_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_5_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_5_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_5_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_5_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_6_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_6_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_6_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_6_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_7_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_7_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_7_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_7_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_8_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_8_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_8_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_8_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_9_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_9_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_9_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_9_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_10_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_10_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_10_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_10_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_11_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_11_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_11_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_11_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_12_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_12_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_12_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_12_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_13_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_13_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_13_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_13_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_14_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_14_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_14_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_14_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_15_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_15_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_15_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_15_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_16_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_16_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_16_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_16_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_17_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_17_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_17_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_17_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_18_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_18_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_18_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_18_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_19_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_19_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_19_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_19_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_20_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_20_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_20_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_20_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_21_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_21_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_21_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_21_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_22_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_22_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_22_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_22_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_23_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_23_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_23_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_23_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_24_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_24_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_24_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_24_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_25_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_25_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_25_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_25_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_26_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_26_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_26_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_26_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_27_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_27_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_27_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_27_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_28_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_28_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_28_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_28_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_29_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_29_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_29_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_29_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_30_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_30_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_30_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_30_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_31_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_31_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_31_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_31_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_32_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_32_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_32_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_32_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_33_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_33_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_33_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_33_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_34_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_34_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_34_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_34_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_35_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_35_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_35_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_35_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_36_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_36_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_36_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_36_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_37_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_37_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_37_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_37_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_38_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_38_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_38_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_38_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_39_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_39_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_39_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_39_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_40_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_40_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_40_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_40_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_41_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_41_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_41_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_41_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_42_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_42_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_42_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_42_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_43_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_43_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_43_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_43_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_44_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_44_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_44_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_44_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_45_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_45_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_45_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_45_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_46_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_46_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_46_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_46_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_47_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_47_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_47_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_47_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_48_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_48_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_48_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_48_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_49_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_49_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_49_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_49_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_50_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_50_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_50_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_50_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_51_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_51_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_51_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_51_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_52_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_52_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_52_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_52_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_53_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_53_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_53_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_53_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_54_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_54_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_54_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_54_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_55_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_55_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_55_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_55_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_56_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_56_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_56_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_56_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_57_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_57_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_57_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_57_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_58_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_58_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_58_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_58_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_59_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_59_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_59_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_59_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_60_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_60_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_60_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_60_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_61_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_61_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_61_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_61_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_62_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_62_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_62_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_62_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_63_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_63_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_63_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_63_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_64_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_64_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_64_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_64_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_65_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_65_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_65_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_65_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_66_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_66_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_66_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_66_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_67_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_67_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_67_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_67_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_68_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_68_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_68_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_68_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_69_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_69_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_69_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_69_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_70_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_70_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_70_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_70_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_71_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_71_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_71_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_71_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_72_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_72_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_72_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_72_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_73_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_73_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_73_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_73_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_74_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_74_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_74_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_74_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_75_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_75_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_75_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_75_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_76_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_76_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_76_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_76_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_77_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_77_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_77_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_77_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_78_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_78_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_78_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_78_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_79_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_79_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_79_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_79_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_80_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_80_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_80_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_80_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_81_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_81_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_81_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_81_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_82_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_82_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_82_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_82_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_83_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_83_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_83_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_83_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_84_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_84_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_84_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_84_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_85_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_85_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_85_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_85_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_86_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_86_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_86_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_86_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_87_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_87_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_87_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_87_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_88_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_88_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_88_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_88_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_89_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_89_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_89_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_89_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_90_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_90_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_90_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_90_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_91_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_91_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_91_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_91_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_92_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_92_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_92_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_92_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_93_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_93_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_93_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_93_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_94_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_94_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_94_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_94_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_95_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_95_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_95_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_95_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_96_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_96_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_96_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_96_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_97_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_97_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_97_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_97_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_98_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_98_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_98_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_98_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_99_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_99_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_99_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_99_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_100_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_100_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_100_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_100_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_101_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_101_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_101_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_101_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_102_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_102_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_102_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_102_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_103_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_103_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_103_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_103_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_104_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_104_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_104_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_104_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_105_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_105_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_105_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_105_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_106_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_106_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_106_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_106_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_107_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_107_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_107_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_107_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_108_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_108_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_108_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_108_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_109_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_109_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_109_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_109_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_110_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_110_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_110_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_110_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_111_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_111_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_111_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_111_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_112_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_112_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_112_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_112_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_113_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_113_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_113_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_113_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_114_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_114_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_114_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_114_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_115_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_115_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_115_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_115_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_116_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_116_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_116_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_116_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_117_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_117_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_117_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_117_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_118_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_118_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_118_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_118_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_119_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_119_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_119_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_119_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_120_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_120_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_120_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_120_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_121_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_121_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_121_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_121_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_122_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_122_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_122_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_122_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_123_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_123_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_123_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_123_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_124_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_124_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_124_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_124_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_125_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_125_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_125_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_125_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_126_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_126_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_126_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_126_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_127_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_127_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_127_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_127_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_128_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_128_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_128_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_128_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_129_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_129_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_129_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_129_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_130_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_130_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_130_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_130_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_131_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_131_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_131_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_131_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_132_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_132_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_132_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_132_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_133_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_133_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_133_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_133_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_134_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_134_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_134_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_134_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_135_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_135_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_135_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_135_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_136_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_136_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_136_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_136_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_137_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_137_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_137_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_137_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_138_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_138_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_138_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_138_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_139_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_139_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_139_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_139_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_140_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_140_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_140_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_140_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_141_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_141_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_141_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_141_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_142_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_142_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_142_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_142_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_143_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_143_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_143_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_143_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_144_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_144_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_144_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_144_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_145_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_145_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_145_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_145_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_146_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_146_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_146_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_146_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_147_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_147_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_147_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_147_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_148_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_148_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_148_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_148_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_149_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_149_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_149_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_149_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_150_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_150_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_150_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_150_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_151_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_151_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_151_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_151_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_152_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_152_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_152_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_152_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_153_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_153_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_153_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_153_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_154_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_154_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_154_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_154_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_155_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_155_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_155_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_155_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_156_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_156_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_156_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_156_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_157_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_157_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_157_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_157_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_158_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_158_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_158_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_158_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_159_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_159_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_159_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_159_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_160_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_160_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_160_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_160_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_161_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_161_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_161_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_161_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_162_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_162_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_162_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_162_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_163_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_163_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_163_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_163_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_164_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_164_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_164_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_164_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_165_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_165_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_165_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_165_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_166_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_166_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_166_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_166_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_167_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_167_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_167_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_167_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_168_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_168_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_168_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_168_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_169_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_169_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_169_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_169_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_170_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_170_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_170_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_170_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_171_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_171_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_171_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_171_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_172_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_172_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_172_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_172_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_173_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_173_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_173_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_173_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_174_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_174_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_174_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_174_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_175_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_175_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_175_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_175_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_176_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_176_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_176_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_176_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_177_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_177_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_177_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_177_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_178_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_178_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_178_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_178_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_179_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_179_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_179_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_179_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_180_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_180_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_180_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_180_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_181_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_181_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_181_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_181_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_182_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_182_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_182_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_182_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_183_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_183_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_183_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_183_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_184_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_184_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_184_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_184_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_185_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_185_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_185_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_185_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_186_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_186_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_186_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_186_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_187_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_187_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_187_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_187_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_188_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_188_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_188_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_188_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_189_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_189_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_189_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_189_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_190_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_190_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_190_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_190_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_191_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_191_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_191_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_191_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_192_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_192_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_192_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_192_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_193_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_193_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_193_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_193_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_194_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_194_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_194_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_194_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_195_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_195_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_195_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_195_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_196_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_196_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_196_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_196_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_197_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_197_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_197_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_197_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_198_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_198_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_198_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_198_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_199_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_199_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_199_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_199_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_200_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_200_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_200_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_200_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_201_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_201_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_201_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_201_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_202_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_202_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_202_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_202_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_203_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_203_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_203_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_203_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_204_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_204_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_204_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_204_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_205_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_205_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_205_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_205_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_206_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_206_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_206_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_206_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_207_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_207_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_207_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_207_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_208_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_208_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_208_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_208_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_209_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_209_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_209_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_209_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_210_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_210_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_210_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_210_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_211_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_211_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_211_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_211_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_212_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_212_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_212_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_212_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_213_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_213_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_213_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_213_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_214_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_214_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_214_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_214_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_215_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_215_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_215_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_215_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_216_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_216_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_216_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_216_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_217_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_217_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_217_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_217_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_218_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_218_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_218_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_218_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_219_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_219_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_219_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_219_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_220_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_220_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_220_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_220_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_221_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_221_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_221_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_221_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_222_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_222_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_222_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_222_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_223_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_223_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_223_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_223_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_224_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_224_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_224_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_224_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_225_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_225_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_225_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_225_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_226_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_226_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_226_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_226_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_227_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_227_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_227_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_227_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_228_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_228_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_228_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_228_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_229_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_229_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_229_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_229_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_230_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_230_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_230_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_230_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_231_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_231_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_231_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_231_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_232_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_232_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_232_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_232_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_233_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_233_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_233_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_233_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_234_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_234_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_234_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_234_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_235_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_235_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_235_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_235_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_236_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_236_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_236_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_236_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_237_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_237_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_237_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_237_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_238_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_238_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_238_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_238_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_239_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_239_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_239_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_239_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_240_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_240_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_240_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_240_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_241_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_241_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_241_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_241_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_242_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_242_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_242_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_242_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_243_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_243_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_243_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_243_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_244_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_244_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_244_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_244_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_245_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_245_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_245_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_245_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_246_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_246_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_246_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_246_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_247_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_247_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_247_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_247_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_248_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_248_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_248_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_248_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_249_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_249_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_249_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_249_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_250_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_250_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_250_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_250_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_251_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_251_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_251_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_251_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_252_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_252_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_252_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_252_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_253_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_253_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_253_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_253_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_254_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_254_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_254_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_254_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_255_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_255_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_255_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_255_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_256_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_256_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_256_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_256_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_257_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_257_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_257_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_257_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_258_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_258_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_258_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_258_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_259_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_259_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_259_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_259_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_260_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_260_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_260_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_260_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_261_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_261_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_261_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_261_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_262_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_262_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_262_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_262_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_263_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_263_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_263_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_263_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_264_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_264_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_264_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_264_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_265_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_265_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_265_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_265_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_266_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_266_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_266_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_266_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_267_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_267_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_267_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_267_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_268_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_268_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_268_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_268_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_269_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_269_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_269_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_269_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_270_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_270_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_270_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_270_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_271_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_271_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_271_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_271_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_272_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_272_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_272_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_272_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_273_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_273_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_273_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_273_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_274_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_274_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_274_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_274_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_275_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_275_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_275_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_275_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_276_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_276_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_276_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_276_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_277_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_277_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_277_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_277_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_278_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_278_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_278_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_278_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_279_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_279_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_279_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_279_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_280_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_280_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_280_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_280_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_281_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_281_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_281_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_281_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_282_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_282_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_282_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_282_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_283_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_283_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_283_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_283_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_284_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_284_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_284_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_284_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_285_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_285_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_285_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_285_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_286_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_286_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_286_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_286_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_287_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_287_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_287_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_287_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_288_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_288_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_288_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_288_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_289_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_289_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_289_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_289_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_290_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_290_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_290_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_290_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_291_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_291_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_291_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_291_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_292_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_292_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_292_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_292_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_293_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_293_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_293_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_293_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_294_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_294_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_294_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_294_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_295_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_295_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_295_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_295_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_296_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_296_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_296_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_296_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_297_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_297_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_297_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_297_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_298_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_298_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_298_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_298_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_299_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_299_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_299_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_299_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_300_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_300_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_300_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_300_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_301_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_301_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_301_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_301_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_302_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_302_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_302_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_302_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_303_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_303_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_303_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_303_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_304_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_304_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_304_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_304_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_305_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_305_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_305_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_305_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_306_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_306_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_306_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_306_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_307_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_307_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_307_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_307_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_308_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_308_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_308_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_308_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_309_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_309_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_309_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_309_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_310_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_310_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_310_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_310_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_311_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_311_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_311_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_311_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_312_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_312_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_312_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_312_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_313_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_313_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_313_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_313_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_314_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_314_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_314_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_314_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_315_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_315_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_315_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_315_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_316_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_316_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_316_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_316_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_317_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_317_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_317_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_317_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_318_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_318_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_318_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_318_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_319_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_319_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_319_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_319_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_320_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_320_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_320_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_320_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_321_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_321_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_321_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_321_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_322_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_322_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_322_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_322_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_323_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_323_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_323_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_323_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_324_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_324_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_324_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_324_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_325_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_325_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_325_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_325_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_326_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_326_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_326_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_326_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_327_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_327_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_327_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_327_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_328_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_328_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_328_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_328_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_329_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_329_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_329_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_329_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_330_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_330_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_330_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_330_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_331_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_331_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_331_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_331_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_332_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_332_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_332_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_332_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_333_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_333_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_333_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_333_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_334_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_334_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_334_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_334_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_335_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_335_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_335_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_335_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_336_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_336_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_336_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_336_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_337_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_337_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_337_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_337_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_338_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_338_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_338_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_338_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_339_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_339_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_339_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_339_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_340_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_340_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_340_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_340_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_341_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_341_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_341_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_341_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_342_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_342_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_342_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_342_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_343_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_343_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_343_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_343_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_344_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_344_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_344_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_344_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_345_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_345_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_345_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_345_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_346_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_346_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_346_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_346_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_347_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_347_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_347_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_347_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_348_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_348_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_348_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_348_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_349_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_349_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_349_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_349_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_350_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_350_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_350_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_350_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_351_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_351_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_351_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_351_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_352_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_352_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_352_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_352_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_353_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_353_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_353_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_353_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_354_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_354_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_354_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_354_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_355_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_355_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_355_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_355_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_356_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_356_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_356_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_356_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_357_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_357_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_357_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_357_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_358_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_358_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_358_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_358_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_359_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_359_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_359_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_359_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_360_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_360_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_360_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_360_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_361_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_361_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_361_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_361_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_362_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_362_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_362_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_362_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_363_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_363_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_363_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_363_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_364_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_364_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_364_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_364_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_365_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_365_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_365_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_365_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_366_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_366_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_366_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_366_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_367_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_367_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_367_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_367_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_368_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_368_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_368_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_368_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_369_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_369_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_369_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_369_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_370_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_370_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_370_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_370_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_371_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_371_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_371_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_371_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_372_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_372_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_372_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_372_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_373_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_373_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_373_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_373_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_374_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_374_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_374_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_374_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_375_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_375_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_375_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_375_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_376_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_376_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_376_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_376_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_377_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_377_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_377_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_377_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_378_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_378_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_378_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_378_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_379_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_379_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_379_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_379_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_380_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_380_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_380_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_380_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_381_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_381_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_381_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_381_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_382_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_382_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_382_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_382_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_383_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_383_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_383_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_383_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_384_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_384_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_384_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_384_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_385_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_385_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_385_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_385_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_386_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_386_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_386_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_386_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_387_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_387_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_387_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_387_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_388_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_388_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_388_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_388_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_389_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_389_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_389_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_389_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_390_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_390_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_390_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_390_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_391_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_391_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_391_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_391_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_392_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_392_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_392_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_392_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_393_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_393_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_393_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_393_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_394_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_394_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_394_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_394_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_395_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_395_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_395_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_395_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_396_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_396_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_396_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_396_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_397_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_397_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_397_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_397_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_398_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_398_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_398_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_398_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_399_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_399_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_399_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_399_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_400_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_400_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_400_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_400_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_401_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_401_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_401_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_401_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_402_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_402_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_402_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_402_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_403_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_403_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_403_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_403_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_404_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_404_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_404_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_404_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_405_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_405_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_405_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_405_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_406_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_406_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_406_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_406_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_407_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_407_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_407_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_407_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_408_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_408_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_408_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_408_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_409_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_409_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_409_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_409_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_410_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_410_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_410_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_410_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_411_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_411_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_411_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_411_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_412_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_412_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_412_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_412_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_413_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_413_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_413_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_413_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_414_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_414_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_414_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_414_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_415_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_415_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_415_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_415_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_416_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_416_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_416_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_416_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_417_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_417_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_417_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_417_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_418_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_418_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_418_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_418_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_419_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_419_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_419_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_419_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_420_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_420_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_420_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_420_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_421_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_421_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_421_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_421_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_422_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_422_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_422_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_422_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_423_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_423_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_423_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_423_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_424_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_424_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_424_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_424_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_425_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_425_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_425_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_425_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_426_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_426_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_426_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_426_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_427_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_427_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_427_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_427_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_428_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_428_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_428_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_428_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_429_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_429_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_429_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_429_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_430_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_430_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_430_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_430_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_431_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_431_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_431_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_431_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_432_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_432_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_432_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_432_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_433_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_433_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_433_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_433_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_434_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_434_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_434_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_434_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_435_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_435_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_435_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_435_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_436_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_436_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_436_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_436_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_437_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_437_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_437_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_437_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_438_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_438_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_438_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_438_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_439_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_439_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_439_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_439_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_440_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_440_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_440_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_440_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_441_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_441_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_441_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_441_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_442_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_442_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_442_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_442_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_443_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_443_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_443_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_443_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_444_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_444_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_444_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_444_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_445_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_445_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_445_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_445_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_446_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_446_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_446_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_446_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_447_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_447_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_447_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_447_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_448_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_448_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_448_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_448_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_449_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_449_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_449_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_449_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_450_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_450_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_450_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_450_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_451_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_451_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_451_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_451_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_452_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_452_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_452_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_452_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_453_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_453_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_453_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_453_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_454_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_454_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_454_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_454_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_455_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_455_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_455_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_455_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_456_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_456_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_456_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_456_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_457_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_457_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_457_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_457_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_458_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_458_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_458_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_458_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_459_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_459_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_459_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_459_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_460_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_460_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_460_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_460_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_461_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_461_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_461_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_461_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_462_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_462_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_462_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_462_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_463_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_463_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_463_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_463_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_464_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_464_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_464_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_464_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_465_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_465_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_465_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_465_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_466_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_466_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_466_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_466_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_467_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_467_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_467_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_467_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_468_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_468_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_468_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_468_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_469_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_469_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_469_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_469_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_470_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_470_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_470_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_470_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_471_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_471_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_471_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_471_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_472_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_472_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_472_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_472_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_473_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_473_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_473_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_473_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_474_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_474_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_474_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_474_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_475_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_475_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_475_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_475_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_476_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_476_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_476_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_476_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_477_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_477_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_477_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_477_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_478_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_478_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_478_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_478_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_479_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_479_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_479_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_479_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_480_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_480_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_480_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_480_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_481_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_481_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_481_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_481_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_482_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_482_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_482_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_482_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_483_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_483_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_483_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_483_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_484_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_484_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_484_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_484_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_485_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_485_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_485_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_485_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_486_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_486_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_486_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_486_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_487_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_487_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_487_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_487_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_488_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_488_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_488_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_488_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_489_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_489_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_489_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_489_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_490_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_490_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_490_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_490_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_491_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_491_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_491_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_491_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_492_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_492_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_492_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_492_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_493_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_493_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_493_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_493_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_494_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_494_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_494_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_494_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_495_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_495_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_495_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_495_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_496_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_496_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_496_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_496_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_497_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_497_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_497_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_497_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_498_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_498_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_498_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_498_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_499_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_499_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_499_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_499_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_500_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_500_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_500_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_500_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_501_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_501_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_501_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_501_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_502_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_502_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_502_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_502_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_503_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_503_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_503_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_503_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_504_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_504_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_504_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_504_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_505_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_505_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_505_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_505_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_506_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_506_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_506_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_506_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_507_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_507_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_507_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_507_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_508_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_508_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_508_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_508_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_509_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_509_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_509_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_509_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_510_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_510_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_510_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_510_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_511_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_511_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_511_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_511_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_512_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_512_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_512_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_512_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_513_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_513_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_513_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_513_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_514_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_514_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_514_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_514_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_515_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_515_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_515_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_515_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_516_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_516_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_516_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_516_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_517_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_517_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_517_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_517_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_518_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_518_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_518_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_518_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_519_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_519_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_519_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_519_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_520_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_520_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_520_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_520_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_521_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_521_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_521_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_521_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_522_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_522_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_522_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_522_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_523_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_523_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_523_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_523_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_524_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_524_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_524_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_524_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_525_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_525_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_525_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_525_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_526_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_526_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_526_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_526_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_527_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_527_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_527_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_527_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_528_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_528_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_528_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_528_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_529_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_529_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_529_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_529_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_530_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_530_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_530_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_530_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_531_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_531_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_531_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_531_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_532_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_532_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_532_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_532_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_533_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_533_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_533_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_533_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_534_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_534_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_534_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_534_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_535_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_535_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_535_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_535_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_536_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_536_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_536_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_536_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_537_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_537_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_537_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_537_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_538_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_538_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_538_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_538_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_539_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_539_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_539_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_539_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_540_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_540_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_540_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_540_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_541_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_541_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_541_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_541_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_542_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_542_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_542_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_542_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_543_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_543_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_543_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_543_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_544_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_544_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_544_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_544_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_545_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_545_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_545_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_545_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_546_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_546_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_546_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_546_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_547_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_547_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_547_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_547_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_548_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_548_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_548_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_548_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_549_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_549_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_549_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_549_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_550_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_550_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_550_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_550_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_551_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_551_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_551_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_551_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_552_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_552_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_552_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_552_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_553_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_553_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_553_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_553_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_554_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_554_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_554_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_554_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_555_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_555_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_555_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_555_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_556_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_556_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_556_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_556_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_557_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_557_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_557_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_557_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_558_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_558_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_558_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_558_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_559_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_559_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_559_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_559_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_560_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_560_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_560_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_560_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_561_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_561_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_561_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_561_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_562_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_562_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_562_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_562_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_563_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_563_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_563_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_563_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_564_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_564_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_564_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_564_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_565_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_565_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_565_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_565_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_566_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_566_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_566_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_566_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_567_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_567_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_567_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_567_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_568_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_568_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_568_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_568_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_569_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_569_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_569_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_569_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_570_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_570_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_570_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_570_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_571_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_571_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_571_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_571_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_572_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_572_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_572_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_572_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_573_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_573_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_573_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_573_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_574_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_574_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_574_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_574_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_575_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_575_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_575_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_575_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_576_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_576_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_576_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_576_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_577_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_577_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_577_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_577_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_578_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_578_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_578_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_578_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_579_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_579_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_579_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_579_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_580_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_580_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_580_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_580_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_581_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_581_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_581_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_581_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_582_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_582_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_582_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_582_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_583_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_583_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_583_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_583_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_584_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_584_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_584_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_584_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_585_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_585_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_585_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_585_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_586_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_586_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_586_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_586_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_587_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_587_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_587_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_587_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_588_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_588_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_588_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_588_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_589_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_589_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_589_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_589_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_590_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_590_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_590_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_590_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_591_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_591_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_591_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_591_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_592_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_592_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_592_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_592_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_593_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_593_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_593_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_593_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_594_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_594_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_594_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_594_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_595_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_595_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_595_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_595_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_596_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_596_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_596_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_596_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_597_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_597_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_597_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_597_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_598_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_598_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_598_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_598_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_599_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_599_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_599_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_599_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_600_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_600_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_600_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_600_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_601_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_601_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_601_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_601_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_602_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_602_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_602_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_602_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_603_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_603_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_603_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_603_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_604_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_604_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_604_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_604_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_605_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_605_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_605_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_605_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_606_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_606_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_606_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_606_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_607_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_607_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_607_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_607_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_608_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_608_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_608_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_608_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_609_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_609_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_609_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_609_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_610_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_610_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_610_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_610_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_611_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_611_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_611_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_611_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_612_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_612_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_612_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_612_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_613_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_613_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_613_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_613_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_614_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_614_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_614_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_614_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_615_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_615_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_615_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_615_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_616_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_616_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_616_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_616_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_617_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_617_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_617_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_617_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_618_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_618_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_618_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_618_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_619_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_619_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_619_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_619_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_620_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_620_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_620_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_620_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_621_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_621_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_621_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_621_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_622_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_622_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_622_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_622_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_623_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_623_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_623_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_623_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_624_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_624_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_624_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_624_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_625_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_625_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_625_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_625_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_626_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_626_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_626_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_626_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_627_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_627_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_627_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_627_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_628_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_628_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_628_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_628_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_629_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_629_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_629_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_629_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_630_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_630_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_630_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_630_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_631_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_631_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_631_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_631_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_632_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_632_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_632_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_632_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_633_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_633_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_633_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_633_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_634_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_634_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_634_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_634_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_635_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_635_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_635_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_635_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_636_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_636_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_636_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_636_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_637_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_637_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_637_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_637_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_638_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_638_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_638_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_638_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_639_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_639_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_639_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_639_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_640_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_640_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_640_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_640_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_641_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_641_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_641_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_641_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_642_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_642_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_642_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_642_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_643_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_643_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_643_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_643_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_644_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_644_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_644_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_644_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_645_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_645_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_645_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_645_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_646_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_646_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_646_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_646_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_647_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_647_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_647_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_647_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_648_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_648_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_648_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_648_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_649_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_649_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_649_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_649_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_650_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_650_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_650_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_650_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_651_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_651_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_651_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_651_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_652_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_652_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_652_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_652_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_653_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_653_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_653_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_653_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_654_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_654_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_654_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_654_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_655_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_655_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_655_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_655_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_656_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_656_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_656_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_656_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_657_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_657_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_657_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_657_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_658_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_658_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_658_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_658_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_659_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_659_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_659_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_659_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_660_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_660_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_660_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_660_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_661_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_661_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_661_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_661_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_662_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_662_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_662_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_662_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_663_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_663_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_663_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_663_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_664_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_664_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_664_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_664_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_665_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_665_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_665_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_665_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_666_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_666_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_666_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_666_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_667_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_667_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_667_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_667_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_668_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_668_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_668_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_668_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_669_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_669_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_669_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_669_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_670_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_670_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_670_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_670_io_z1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_671_io_a0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_671_io_a1; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_671_io_z0; // @[bitonic_sort.scala 31:25]
  wire [7:0] Swapper_671_io_z1; // @[bitonic_sort.scala 31:25]
  Swapper Swapper ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_io_a0),
    .io_a1(Swapper_io_a1),
    .io_z0(Swapper_io_z0),
    .io_z1(Swapper_io_z1)
  );
  Swapper Swapper_1 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_1_io_a0),
    .io_a1(Swapper_1_io_a1),
    .io_z0(Swapper_1_io_z0),
    .io_z1(Swapper_1_io_z1)
  );
  Swapper Swapper_2 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_2_io_a0),
    .io_a1(Swapper_2_io_a1),
    .io_z0(Swapper_2_io_z0),
    .io_z1(Swapper_2_io_z1)
  );
  Swapper Swapper_3 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_3_io_a0),
    .io_a1(Swapper_3_io_a1),
    .io_z0(Swapper_3_io_z0),
    .io_z1(Swapper_3_io_z1)
  );
  Swapper Swapper_4 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_4_io_a0),
    .io_a1(Swapper_4_io_a1),
    .io_z0(Swapper_4_io_z0),
    .io_z1(Swapper_4_io_z1)
  );
  Swapper Swapper_5 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_5_io_a0),
    .io_a1(Swapper_5_io_a1),
    .io_z0(Swapper_5_io_z0),
    .io_z1(Swapper_5_io_z1)
  );
  Swapper Swapper_6 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_6_io_a0),
    .io_a1(Swapper_6_io_a1),
    .io_z0(Swapper_6_io_z0),
    .io_z1(Swapper_6_io_z1)
  );
  Swapper Swapper_7 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_7_io_a0),
    .io_a1(Swapper_7_io_a1),
    .io_z0(Swapper_7_io_z0),
    .io_z1(Swapper_7_io_z1)
  );
  Swapper Swapper_8 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_8_io_a0),
    .io_a1(Swapper_8_io_a1),
    .io_z0(Swapper_8_io_z0),
    .io_z1(Swapper_8_io_z1)
  );
  Swapper Swapper_9 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_9_io_a0),
    .io_a1(Swapper_9_io_a1),
    .io_z0(Swapper_9_io_z0),
    .io_z1(Swapper_9_io_z1)
  );
  Swapper Swapper_10 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_10_io_a0),
    .io_a1(Swapper_10_io_a1),
    .io_z0(Swapper_10_io_z0),
    .io_z1(Swapper_10_io_z1)
  );
  Swapper Swapper_11 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_11_io_a0),
    .io_a1(Swapper_11_io_a1),
    .io_z0(Swapper_11_io_z0),
    .io_z1(Swapper_11_io_z1)
  );
  Swapper Swapper_12 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_12_io_a0),
    .io_a1(Swapper_12_io_a1),
    .io_z0(Swapper_12_io_z0),
    .io_z1(Swapper_12_io_z1)
  );
  Swapper Swapper_13 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_13_io_a0),
    .io_a1(Swapper_13_io_a1),
    .io_z0(Swapper_13_io_z0),
    .io_z1(Swapper_13_io_z1)
  );
  Swapper Swapper_14 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_14_io_a0),
    .io_a1(Swapper_14_io_a1),
    .io_z0(Swapper_14_io_z0),
    .io_z1(Swapper_14_io_z1)
  );
  Swapper Swapper_15 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_15_io_a0),
    .io_a1(Swapper_15_io_a1),
    .io_z0(Swapper_15_io_z0),
    .io_z1(Swapper_15_io_z1)
  );
  Swapper Swapper_16 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_16_io_a0),
    .io_a1(Swapper_16_io_a1),
    .io_z0(Swapper_16_io_z0),
    .io_z1(Swapper_16_io_z1)
  );
  Swapper Swapper_17 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_17_io_a0),
    .io_a1(Swapper_17_io_a1),
    .io_z0(Swapper_17_io_z0),
    .io_z1(Swapper_17_io_z1)
  );
  Swapper Swapper_18 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_18_io_a0),
    .io_a1(Swapper_18_io_a1),
    .io_z0(Swapper_18_io_z0),
    .io_z1(Swapper_18_io_z1)
  );
  Swapper Swapper_19 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_19_io_a0),
    .io_a1(Swapper_19_io_a1),
    .io_z0(Swapper_19_io_z0),
    .io_z1(Swapper_19_io_z1)
  );
  Swapper Swapper_20 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_20_io_a0),
    .io_a1(Swapper_20_io_a1),
    .io_z0(Swapper_20_io_z0),
    .io_z1(Swapper_20_io_z1)
  );
  Swapper Swapper_21 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_21_io_a0),
    .io_a1(Swapper_21_io_a1),
    .io_z0(Swapper_21_io_z0),
    .io_z1(Swapper_21_io_z1)
  );
  Swapper Swapper_22 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_22_io_a0),
    .io_a1(Swapper_22_io_a1),
    .io_z0(Swapper_22_io_z0),
    .io_z1(Swapper_22_io_z1)
  );
  Swapper Swapper_23 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_23_io_a0),
    .io_a1(Swapper_23_io_a1),
    .io_z0(Swapper_23_io_z0),
    .io_z1(Swapper_23_io_z1)
  );
  Swapper Swapper_24 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_24_io_a0),
    .io_a1(Swapper_24_io_a1),
    .io_z0(Swapper_24_io_z0),
    .io_z1(Swapper_24_io_z1)
  );
  Swapper Swapper_25 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_25_io_a0),
    .io_a1(Swapper_25_io_a1),
    .io_z0(Swapper_25_io_z0),
    .io_z1(Swapper_25_io_z1)
  );
  Swapper Swapper_26 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_26_io_a0),
    .io_a1(Swapper_26_io_a1),
    .io_z0(Swapper_26_io_z0),
    .io_z1(Swapper_26_io_z1)
  );
  Swapper Swapper_27 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_27_io_a0),
    .io_a1(Swapper_27_io_a1),
    .io_z0(Swapper_27_io_z0),
    .io_z1(Swapper_27_io_z1)
  );
  Swapper Swapper_28 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_28_io_a0),
    .io_a1(Swapper_28_io_a1),
    .io_z0(Swapper_28_io_z0),
    .io_z1(Swapper_28_io_z1)
  );
  Swapper Swapper_29 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_29_io_a0),
    .io_a1(Swapper_29_io_a1),
    .io_z0(Swapper_29_io_z0),
    .io_z1(Swapper_29_io_z1)
  );
  Swapper Swapper_30 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_30_io_a0),
    .io_a1(Swapper_30_io_a1),
    .io_z0(Swapper_30_io_z0),
    .io_z1(Swapper_30_io_z1)
  );
  Swapper Swapper_31 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_31_io_a0),
    .io_a1(Swapper_31_io_a1),
    .io_z0(Swapper_31_io_z0),
    .io_z1(Swapper_31_io_z1)
  );
  Swapper Swapper_32 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_32_io_a0),
    .io_a1(Swapper_32_io_a1),
    .io_z0(Swapper_32_io_z0),
    .io_z1(Swapper_32_io_z1)
  );
  Swapper Swapper_33 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_33_io_a0),
    .io_a1(Swapper_33_io_a1),
    .io_z0(Swapper_33_io_z0),
    .io_z1(Swapper_33_io_z1)
  );
  Swapper Swapper_34 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_34_io_a0),
    .io_a1(Swapper_34_io_a1),
    .io_z0(Swapper_34_io_z0),
    .io_z1(Swapper_34_io_z1)
  );
  Swapper Swapper_35 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_35_io_a0),
    .io_a1(Swapper_35_io_a1),
    .io_z0(Swapper_35_io_z0),
    .io_z1(Swapper_35_io_z1)
  );
  Swapper Swapper_36 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_36_io_a0),
    .io_a1(Swapper_36_io_a1),
    .io_z0(Swapper_36_io_z0),
    .io_z1(Swapper_36_io_z1)
  );
  Swapper Swapper_37 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_37_io_a0),
    .io_a1(Swapper_37_io_a1),
    .io_z0(Swapper_37_io_z0),
    .io_z1(Swapper_37_io_z1)
  );
  Swapper Swapper_38 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_38_io_a0),
    .io_a1(Swapper_38_io_a1),
    .io_z0(Swapper_38_io_z0),
    .io_z1(Swapper_38_io_z1)
  );
  Swapper Swapper_39 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_39_io_a0),
    .io_a1(Swapper_39_io_a1),
    .io_z0(Swapper_39_io_z0),
    .io_z1(Swapper_39_io_z1)
  );
  Swapper Swapper_40 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_40_io_a0),
    .io_a1(Swapper_40_io_a1),
    .io_z0(Swapper_40_io_z0),
    .io_z1(Swapper_40_io_z1)
  );
  Swapper Swapper_41 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_41_io_a0),
    .io_a1(Swapper_41_io_a1),
    .io_z0(Swapper_41_io_z0),
    .io_z1(Swapper_41_io_z1)
  );
  Swapper Swapper_42 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_42_io_a0),
    .io_a1(Swapper_42_io_a1),
    .io_z0(Swapper_42_io_z0),
    .io_z1(Swapper_42_io_z1)
  );
  Swapper Swapper_43 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_43_io_a0),
    .io_a1(Swapper_43_io_a1),
    .io_z0(Swapper_43_io_z0),
    .io_z1(Swapper_43_io_z1)
  );
  Swapper Swapper_44 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_44_io_a0),
    .io_a1(Swapper_44_io_a1),
    .io_z0(Swapper_44_io_z0),
    .io_z1(Swapper_44_io_z1)
  );
  Swapper Swapper_45 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_45_io_a0),
    .io_a1(Swapper_45_io_a1),
    .io_z0(Swapper_45_io_z0),
    .io_z1(Swapper_45_io_z1)
  );
  Swapper Swapper_46 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_46_io_a0),
    .io_a1(Swapper_46_io_a1),
    .io_z0(Swapper_46_io_z0),
    .io_z1(Swapper_46_io_z1)
  );
  Swapper Swapper_47 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_47_io_a0),
    .io_a1(Swapper_47_io_a1),
    .io_z0(Swapper_47_io_z0),
    .io_z1(Swapper_47_io_z1)
  );
  Swapper Swapper_48 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_48_io_a0),
    .io_a1(Swapper_48_io_a1),
    .io_z0(Swapper_48_io_z0),
    .io_z1(Swapper_48_io_z1)
  );
  Swapper Swapper_49 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_49_io_a0),
    .io_a1(Swapper_49_io_a1),
    .io_z0(Swapper_49_io_z0),
    .io_z1(Swapper_49_io_z1)
  );
  Swapper Swapper_50 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_50_io_a0),
    .io_a1(Swapper_50_io_a1),
    .io_z0(Swapper_50_io_z0),
    .io_z1(Swapper_50_io_z1)
  );
  Swapper Swapper_51 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_51_io_a0),
    .io_a1(Swapper_51_io_a1),
    .io_z0(Swapper_51_io_z0),
    .io_z1(Swapper_51_io_z1)
  );
  Swapper Swapper_52 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_52_io_a0),
    .io_a1(Swapper_52_io_a1),
    .io_z0(Swapper_52_io_z0),
    .io_z1(Swapper_52_io_z1)
  );
  Swapper Swapper_53 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_53_io_a0),
    .io_a1(Swapper_53_io_a1),
    .io_z0(Swapper_53_io_z0),
    .io_z1(Swapper_53_io_z1)
  );
  Swapper Swapper_54 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_54_io_a0),
    .io_a1(Swapper_54_io_a1),
    .io_z0(Swapper_54_io_z0),
    .io_z1(Swapper_54_io_z1)
  );
  Swapper Swapper_55 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_55_io_a0),
    .io_a1(Swapper_55_io_a1),
    .io_z0(Swapper_55_io_z0),
    .io_z1(Swapper_55_io_z1)
  );
  Swapper Swapper_56 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_56_io_a0),
    .io_a1(Swapper_56_io_a1),
    .io_z0(Swapper_56_io_z0),
    .io_z1(Swapper_56_io_z1)
  );
  Swapper Swapper_57 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_57_io_a0),
    .io_a1(Swapper_57_io_a1),
    .io_z0(Swapper_57_io_z0),
    .io_z1(Swapper_57_io_z1)
  );
  Swapper Swapper_58 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_58_io_a0),
    .io_a1(Swapper_58_io_a1),
    .io_z0(Swapper_58_io_z0),
    .io_z1(Swapper_58_io_z1)
  );
  Swapper Swapper_59 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_59_io_a0),
    .io_a1(Swapper_59_io_a1),
    .io_z0(Swapper_59_io_z0),
    .io_z1(Swapper_59_io_z1)
  );
  Swapper Swapper_60 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_60_io_a0),
    .io_a1(Swapper_60_io_a1),
    .io_z0(Swapper_60_io_z0),
    .io_z1(Swapper_60_io_z1)
  );
  Swapper Swapper_61 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_61_io_a0),
    .io_a1(Swapper_61_io_a1),
    .io_z0(Swapper_61_io_z0),
    .io_z1(Swapper_61_io_z1)
  );
  Swapper Swapper_62 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_62_io_a0),
    .io_a1(Swapper_62_io_a1),
    .io_z0(Swapper_62_io_z0),
    .io_z1(Swapper_62_io_z1)
  );
  Swapper Swapper_63 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_63_io_a0),
    .io_a1(Swapper_63_io_a1),
    .io_z0(Swapper_63_io_z0),
    .io_z1(Swapper_63_io_z1)
  );
  Swapper Swapper_64 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_64_io_a0),
    .io_a1(Swapper_64_io_a1),
    .io_z0(Swapper_64_io_z0),
    .io_z1(Swapper_64_io_z1)
  );
  Swapper Swapper_65 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_65_io_a0),
    .io_a1(Swapper_65_io_a1),
    .io_z0(Swapper_65_io_z0),
    .io_z1(Swapper_65_io_z1)
  );
  Swapper Swapper_66 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_66_io_a0),
    .io_a1(Swapper_66_io_a1),
    .io_z0(Swapper_66_io_z0),
    .io_z1(Swapper_66_io_z1)
  );
  Swapper Swapper_67 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_67_io_a0),
    .io_a1(Swapper_67_io_a1),
    .io_z0(Swapper_67_io_z0),
    .io_z1(Swapper_67_io_z1)
  );
  Swapper Swapper_68 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_68_io_a0),
    .io_a1(Swapper_68_io_a1),
    .io_z0(Swapper_68_io_z0),
    .io_z1(Swapper_68_io_z1)
  );
  Swapper Swapper_69 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_69_io_a0),
    .io_a1(Swapper_69_io_a1),
    .io_z0(Swapper_69_io_z0),
    .io_z1(Swapper_69_io_z1)
  );
  Swapper Swapper_70 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_70_io_a0),
    .io_a1(Swapper_70_io_a1),
    .io_z0(Swapper_70_io_z0),
    .io_z1(Swapper_70_io_z1)
  );
  Swapper Swapper_71 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_71_io_a0),
    .io_a1(Swapper_71_io_a1),
    .io_z0(Swapper_71_io_z0),
    .io_z1(Swapper_71_io_z1)
  );
  Swapper Swapper_72 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_72_io_a0),
    .io_a1(Swapper_72_io_a1),
    .io_z0(Swapper_72_io_z0),
    .io_z1(Swapper_72_io_z1)
  );
  Swapper Swapper_73 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_73_io_a0),
    .io_a1(Swapper_73_io_a1),
    .io_z0(Swapper_73_io_z0),
    .io_z1(Swapper_73_io_z1)
  );
  Swapper Swapper_74 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_74_io_a0),
    .io_a1(Swapper_74_io_a1),
    .io_z0(Swapper_74_io_z0),
    .io_z1(Swapper_74_io_z1)
  );
  Swapper Swapper_75 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_75_io_a0),
    .io_a1(Swapper_75_io_a1),
    .io_z0(Swapper_75_io_z0),
    .io_z1(Swapper_75_io_z1)
  );
  Swapper Swapper_76 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_76_io_a0),
    .io_a1(Swapper_76_io_a1),
    .io_z0(Swapper_76_io_z0),
    .io_z1(Swapper_76_io_z1)
  );
  Swapper Swapper_77 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_77_io_a0),
    .io_a1(Swapper_77_io_a1),
    .io_z0(Swapper_77_io_z0),
    .io_z1(Swapper_77_io_z1)
  );
  Swapper Swapper_78 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_78_io_a0),
    .io_a1(Swapper_78_io_a1),
    .io_z0(Swapper_78_io_z0),
    .io_z1(Swapper_78_io_z1)
  );
  Swapper Swapper_79 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_79_io_a0),
    .io_a1(Swapper_79_io_a1),
    .io_z0(Swapper_79_io_z0),
    .io_z1(Swapper_79_io_z1)
  );
  Swapper Swapper_80 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_80_io_a0),
    .io_a1(Swapper_80_io_a1),
    .io_z0(Swapper_80_io_z0),
    .io_z1(Swapper_80_io_z1)
  );
  Swapper Swapper_81 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_81_io_a0),
    .io_a1(Swapper_81_io_a1),
    .io_z0(Swapper_81_io_z0),
    .io_z1(Swapper_81_io_z1)
  );
  Swapper Swapper_82 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_82_io_a0),
    .io_a1(Swapper_82_io_a1),
    .io_z0(Swapper_82_io_z0),
    .io_z1(Swapper_82_io_z1)
  );
  Swapper Swapper_83 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_83_io_a0),
    .io_a1(Swapper_83_io_a1),
    .io_z0(Swapper_83_io_z0),
    .io_z1(Swapper_83_io_z1)
  );
  Swapper Swapper_84 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_84_io_a0),
    .io_a1(Swapper_84_io_a1),
    .io_z0(Swapper_84_io_z0),
    .io_z1(Swapper_84_io_z1)
  );
  Swapper Swapper_85 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_85_io_a0),
    .io_a1(Swapper_85_io_a1),
    .io_z0(Swapper_85_io_z0),
    .io_z1(Swapper_85_io_z1)
  );
  Swapper Swapper_86 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_86_io_a0),
    .io_a1(Swapper_86_io_a1),
    .io_z0(Swapper_86_io_z0),
    .io_z1(Swapper_86_io_z1)
  );
  Swapper Swapper_87 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_87_io_a0),
    .io_a1(Swapper_87_io_a1),
    .io_z0(Swapper_87_io_z0),
    .io_z1(Swapper_87_io_z1)
  );
  Swapper Swapper_88 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_88_io_a0),
    .io_a1(Swapper_88_io_a1),
    .io_z0(Swapper_88_io_z0),
    .io_z1(Swapper_88_io_z1)
  );
  Swapper Swapper_89 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_89_io_a0),
    .io_a1(Swapper_89_io_a1),
    .io_z0(Swapper_89_io_z0),
    .io_z1(Swapper_89_io_z1)
  );
  Swapper Swapper_90 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_90_io_a0),
    .io_a1(Swapper_90_io_a1),
    .io_z0(Swapper_90_io_z0),
    .io_z1(Swapper_90_io_z1)
  );
  Swapper Swapper_91 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_91_io_a0),
    .io_a1(Swapper_91_io_a1),
    .io_z0(Swapper_91_io_z0),
    .io_z1(Swapper_91_io_z1)
  );
  Swapper Swapper_92 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_92_io_a0),
    .io_a1(Swapper_92_io_a1),
    .io_z0(Swapper_92_io_z0),
    .io_z1(Swapper_92_io_z1)
  );
  Swapper Swapper_93 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_93_io_a0),
    .io_a1(Swapper_93_io_a1),
    .io_z0(Swapper_93_io_z0),
    .io_z1(Swapper_93_io_z1)
  );
  Swapper Swapper_94 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_94_io_a0),
    .io_a1(Swapper_94_io_a1),
    .io_z0(Swapper_94_io_z0),
    .io_z1(Swapper_94_io_z1)
  );
  Swapper Swapper_95 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_95_io_a0),
    .io_a1(Swapper_95_io_a1),
    .io_z0(Swapper_95_io_z0),
    .io_z1(Swapper_95_io_z1)
  );
  Swapper Swapper_96 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_96_io_a0),
    .io_a1(Swapper_96_io_a1),
    .io_z0(Swapper_96_io_z0),
    .io_z1(Swapper_96_io_z1)
  );
  Swapper Swapper_97 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_97_io_a0),
    .io_a1(Swapper_97_io_a1),
    .io_z0(Swapper_97_io_z0),
    .io_z1(Swapper_97_io_z1)
  );
  Swapper Swapper_98 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_98_io_a0),
    .io_a1(Swapper_98_io_a1),
    .io_z0(Swapper_98_io_z0),
    .io_z1(Swapper_98_io_z1)
  );
  Swapper Swapper_99 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_99_io_a0),
    .io_a1(Swapper_99_io_a1),
    .io_z0(Swapper_99_io_z0),
    .io_z1(Swapper_99_io_z1)
  );
  Swapper Swapper_100 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_100_io_a0),
    .io_a1(Swapper_100_io_a1),
    .io_z0(Swapper_100_io_z0),
    .io_z1(Swapper_100_io_z1)
  );
  Swapper Swapper_101 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_101_io_a0),
    .io_a1(Swapper_101_io_a1),
    .io_z0(Swapper_101_io_z0),
    .io_z1(Swapper_101_io_z1)
  );
  Swapper Swapper_102 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_102_io_a0),
    .io_a1(Swapper_102_io_a1),
    .io_z0(Swapper_102_io_z0),
    .io_z1(Swapper_102_io_z1)
  );
  Swapper Swapper_103 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_103_io_a0),
    .io_a1(Swapper_103_io_a1),
    .io_z0(Swapper_103_io_z0),
    .io_z1(Swapper_103_io_z1)
  );
  Swapper Swapper_104 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_104_io_a0),
    .io_a1(Swapper_104_io_a1),
    .io_z0(Swapper_104_io_z0),
    .io_z1(Swapper_104_io_z1)
  );
  Swapper Swapper_105 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_105_io_a0),
    .io_a1(Swapper_105_io_a1),
    .io_z0(Swapper_105_io_z0),
    .io_z1(Swapper_105_io_z1)
  );
  Swapper Swapper_106 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_106_io_a0),
    .io_a1(Swapper_106_io_a1),
    .io_z0(Swapper_106_io_z0),
    .io_z1(Swapper_106_io_z1)
  );
  Swapper Swapper_107 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_107_io_a0),
    .io_a1(Swapper_107_io_a1),
    .io_z0(Swapper_107_io_z0),
    .io_z1(Swapper_107_io_z1)
  );
  Swapper Swapper_108 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_108_io_a0),
    .io_a1(Swapper_108_io_a1),
    .io_z0(Swapper_108_io_z0),
    .io_z1(Swapper_108_io_z1)
  );
  Swapper Swapper_109 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_109_io_a0),
    .io_a1(Swapper_109_io_a1),
    .io_z0(Swapper_109_io_z0),
    .io_z1(Swapper_109_io_z1)
  );
  Swapper Swapper_110 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_110_io_a0),
    .io_a1(Swapper_110_io_a1),
    .io_z0(Swapper_110_io_z0),
    .io_z1(Swapper_110_io_z1)
  );
  Swapper Swapper_111 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_111_io_a0),
    .io_a1(Swapper_111_io_a1),
    .io_z0(Swapper_111_io_z0),
    .io_z1(Swapper_111_io_z1)
  );
  Swapper Swapper_112 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_112_io_a0),
    .io_a1(Swapper_112_io_a1),
    .io_z0(Swapper_112_io_z0),
    .io_z1(Swapper_112_io_z1)
  );
  Swapper Swapper_113 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_113_io_a0),
    .io_a1(Swapper_113_io_a1),
    .io_z0(Swapper_113_io_z0),
    .io_z1(Swapper_113_io_z1)
  );
  Swapper Swapper_114 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_114_io_a0),
    .io_a1(Swapper_114_io_a1),
    .io_z0(Swapper_114_io_z0),
    .io_z1(Swapper_114_io_z1)
  );
  Swapper Swapper_115 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_115_io_a0),
    .io_a1(Swapper_115_io_a1),
    .io_z0(Swapper_115_io_z0),
    .io_z1(Swapper_115_io_z1)
  );
  Swapper Swapper_116 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_116_io_a0),
    .io_a1(Swapper_116_io_a1),
    .io_z0(Swapper_116_io_z0),
    .io_z1(Swapper_116_io_z1)
  );
  Swapper Swapper_117 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_117_io_a0),
    .io_a1(Swapper_117_io_a1),
    .io_z0(Swapper_117_io_z0),
    .io_z1(Swapper_117_io_z1)
  );
  Swapper Swapper_118 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_118_io_a0),
    .io_a1(Swapper_118_io_a1),
    .io_z0(Swapper_118_io_z0),
    .io_z1(Swapper_118_io_z1)
  );
  Swapper Swapper_119 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_119_io_a0),
    .io_a1(Swapper_119_io_a1),
    .io_z0(Swapper_119_io_z0),
    .io_z1(Swapper_119_io_z1)
  );
  Swapper Swapper_120 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_120_io_a0),
    .io_a1(Swapper_120_io_a1),
    .io_z0(Swapper_120_io_z0),
    .io_z1(Swapper_120_io_z1)
  );
  Swapper Swapper_121 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_121_io_a0),
    .io_a1(Swapper_121_io_a1),
    .io_z0(Swapper_121_io_z0),
    .io_z1(Swapper_121_io_z1)
  );
  Swapper Swapper_122 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_122_io_a0),
    .io_a1(Swapper_122_io_a1),
    .io_z0(Swapper_122_io_z0),
    .io_z1(Swapper_122_io_z1)
  );
  Swapper Swapper_123 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_123_io_a0),
    .io_a1(Swapper_123_io_a1),
    .io_z0(Swapper_123_io_z0),
    .io_z1(Swapper_123_io_z1)
  );
  Swapper Swapper_124 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_124_io_a0),
    .io_a1(Swapper_124_io_a1),
    .io_z0(Swapper_124_io_z0),
    .io_z1(Swapper_124_io_z1)
  );
  Swapper Swapper_125 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_125_io_a0),
    .io_a1(Swapper_125_io_a1),
    .io_z0(Swapper_125_io_z0),
    .io_z1(Swapper_125_io_z1)
  );
  Swapper Swapper_126 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_126_io_a0),
    .io_a1(Swapper_126_io_a1),
    .io_z0(Swapper_126_io_z0),
    .io_z1(Swapper_126_io_z1)
  );
  Swapper Swapper_127 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_127_io_a0),
    .io_a1(Swapper_127_io_a1),
    .io_z0(Swapper_127_io_z0),
    .io_z1(Swapper_127_io_z1)
  );
  Swapper Swapper_128 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_128_io_a0),
    .io_a1(Swapper_128_io_a1),
    .io_z0(Swapper_128_io_z0),
    .io_z1(Swapper_128_io_z1)
  );
  Swapper Swapper_129 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_129_io_a0),
    .io_a1(Swapper_129_io_a1),
    .io_z0(Swapper_129_io_z0),
    .io_z1(Swapper_129_io_z1)
  );
  Swapper Swapper_130 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_130_io_a0),
    .io_a1(Swapper_130_io_a1),
    .io_z0(Swapper_130_io_z0),
    .io_z1(Swapper_130_io_z1)
  );
  Swapper Swapper_131 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_131_io_a0),
    .io_a1(Swapper_131_io_a1),
    .io_z0(Swapper_131_io_z0),
    .io_z1(Swapper_131_io_z1)
  );
  Swapper Swapper_132 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_132_io_a0),
    .io_a1(Swapper_132_io_a1),
    .io_z0(Swapper_132_io_z0),
    .io_z1(Swapper_132_io_z1)
  );
  Swapper Swapper_133 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_133_io_a0),
    .io_a1(Swapper_133_io_a1),
    .io_z0(Swapper_133_io_z0),
    .io_z1(Swapper_133_io_z1)
  );
  Swapper Swapper_134 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_134_io_a0),
    .io_a1(Swapper_134_io_a1),
    .io_z0(Swapper_134_io_z0),
    .io_z1(Swapper_134_io_z1)
  );
  Swapper Swapper_135 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_135_io_a0),
    .io_a1(Swapper_135_io_a1),
    .io_z0(Swapper_135_io_z0),
    .io_z1(Swapper_135_io_z1)
  );
  Swapper Swapper_136 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_136_io_a0),
    .io_a1(Swapper_136_io_a1),
    .io_z0(Swapper_136_io_z0),
    .io_z1(Swapper_136_io_z1)
  );
  Swapper Swapper_137 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_137_io_a0),
    .io_a1(Swapper_137_io_a1),
    .io_z0(Swapper_137_io_z0),
    .io_z1(Swapper_137_io_z1)
  );
  Swapper Swapper_138 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_138_io_a0),
    .io_a1(Swapper_138_io_a1),
    .io_z0(Swapper_138_io_z0),
    .io_z1(Swapper_138_io_z1)
  );
  Swapper Swapper_139 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_139_io_a0),
    .io_a1(Swapper_139_io_a1),
    .io_z0(Swapper_139_io_z0),
    .io_z1(Swapper_139_io_z1)
  );
  Swapper Swapper_140 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_140_io_a0),
    .io_a1(Swapper_140_io_a1),
    .io_z0(Swapper_140_io_z0),
    .io_z1(Swapper_140_io_z1)
  );
  Swapper Swapper_141 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_141_io_a0),
    .io_a1(Swapper_141_io_a1),
    .io_z0(Swapper_141_io_z0),
    .io_z1(Swapper_141_io_z1)
  );
  Swapper Swapper_142 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_142_io_a0),
    .io_a1(Swapper_142_io_a1),
    .io_z0(Swapper_142_io_z0),
    .io_z1(Swapper_142_io_z1)
  );
  Swapper Swapper_143 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_143_io_a0),
    .io_a1(Swapper_143_io_a1),
    .io_z0(Swapper_143_io_z0),
    .io_z1(Swapper_143_io_z1)
  );
  Swapper Swapper_144 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_144_io_a0),
    .io_a1(Swapper_144_io_a1),
    .io_z0(Swapper_144_io_z0),
    .io_z1(Swapper_144_io_z1)
  );
  Swapper Swapper_145 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_145_io_a0),
    .io_a1(Swapper_145_io_a1),
    .io_z0(Swapper_145_io_z0),
    .io_z1(Swapper_145_io_z1)
  );
  Swapper Swapper_146 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_146_io_a0),
    .io_a1(Swapper_146_io_a1),
    .io_z0(Swapper_146_io_z0),
    .io_z1(Swapper_146_io_z1)
  );
  Swapper Swapper_147 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_147_io_a0),
    .io_a1(Swapper_147_io_a1),
    .io_z0(Swapper_147_io_z0),
    .io_z1(Swapper_147_io_z1)
  );
  Swapper Swapper_148 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_148_io_a0),
    .io_a1(Swapper_148_io_a1),
    .io_z0(Swapper_148_io_z0),
    .io_z1(Swapper_148_io_z1)
  );
  Swapper Swapper_149 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_149_io_a0),
    .io_a1(Swapper_149_io_a1),
    .io_z0(Swapper_149_io_z0),
    .io_z1(Swapper_149_io_z1)
  );
  Swapper Swapper_150 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_150_io_a0),
    .io_a1(Swapper_150_io_a1),
    .io_z0(Swapper_150_io_z0),
    .io_z1(Swapper_150_io_z1)
  );
  Swapper Swapper_151 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_151_io_a0),
    .io_a1(Swapper_151_io_a1),
    .io_z0(Swapper_151_io_z0),
    .io_z1(Swapper_151_io_z1)
  );
  Swapper Swapper_152 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_152_io_a0),
    .io_a1(Swapper_152_io_a1),
    .io_z0(Swapper_152_io_z0),
    .io_z1(Swapper_152_io_z1)
  );
  Swapper Swapper_153 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_153_io_a0),
    .io_a1(Swapper_153_io_a1),
    .io_z0(Swapper_153_io_z0),
    .io_z1(Swapper_153_io_z1)
  );
  Swapper Swapper_154 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_154_io_a0),
    .io_a1(Swapper_154_io_a1),
    .io_z0(Swapper_154_io_z0),
    .io_z1(Swapper_154_io_z1)
  );
  Swapper Swapper_155 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_155_io_a0),
    .io_a1(Swapper_155_io_a1),
    .io_z0(Swapper_155_io_z0),
    .io_z1(Swapper_155_io_z1)
  );
  Swapper Swapper_156 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_156_io_a0),
    .io_a1(Swapper_156_io_a1),
    .io_z0(Swapper_156_io_z0),
    .io_z1(Swapper_156_io_z1)
  );
  Swapper Swapper_157 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_157_io_a0),
    .io_a1(Swapper_157_io_a1),
    .io_z0(Swapper_157_io_z0),
    .io_z1(Swapper_157_io_z1)
  );
  Swapper Swapper_158 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_158_io_a0),
    .io_a1(Swapper_158_io_a1),
    .io_z0(Swapper_158_io_z0),
    .io_z1(Swapper_158_io_z1)
  );
  Swapper Swapper_159 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_159_io_a0),
    .io_a1(Swapper_159_io_a1),
    .io_z0(Swapper_159_io_z0),
    .io_z1(Swapper_159_io_z1)
  );
  Swapper Swapper_160 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_160_io_a0),
    .io_a1(Swapper_160_io_a1),
    .io_z0(Swapper_160_io_z0),
    .io_z1(Swapper_160_io_z1)
  );
  Swapper Swapper_161 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_161_io_a0),
    .io_a1(Swapper_161_io_a1),
    .io_z0(Swapper_161_io_z0),
    .io_z1(Swapper_161_io_z1)
  );
  Swapper Swapper_162 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_162_io_a0),
    .io_a1(Swapper_162_io_a1),
    .io_z0(Swapper_162_io_z0),
    .io_z1(Swapper_162_io_z1)
  );
  Swapper Swapper_163 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_163_io_a0),
    .io_a1(Swapper_163_io_a1),
    .io_z0(Swapper_163_io_z0),
    .io_z1(Swapper_163_io_z1)
  );
  Swapper Swapper_164 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_164_io_a0),
    .io_a1(Swapper_164_io_a1),
    .io_z0(Swapper_164_io_z0),
    .io_z1(Swapper_164_io_z1)
  );
  Swapper Swapper_165 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_165_io_a0),
    .io_a1(Swapper_165_io_a1),
    .io_z0(Swapper_165_io_z0),
    .io_z1(Swapper_165_io_z1)
  );
  Swapper Swapper_166 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_166_io_a0),
    .io_a1(Swapper_166_io_a1),
    .io_z0(Swapper_166_io_z0),
    .io_z1(Swapper_166_io_z1)
  );
  Swapper Swapper_167 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_167_io_a0),
    .io_a1(Swapper_167_io_a1),
    .io_z0(Swapper_167_io_z0),
    .io_z1(Swapper_167_io_z1)
  );
  Swapper Swapper_168 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_168_io_a0),
    .io_a1(Swapper_168_io_a1),
    .io_z0(Swapper_168_io_z0),
    .io_z1(Swapper_168_io_z1)
  );
  Swapper Swapper_169 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_169_io_a0),
    .io_a1(Swapper_169_io_a1),
    .io_z0(Swapper_169_io_z0),
    .io_z1(Swapper_169_io_z1)
  );
  Swapper Swapper_170 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_170_io_a0),
    .io_a1(Swapper_170_io_a1),
    .io_z0(Swapper_170_io_z0),
    .io_z1(Swapper_170_io_z1)
  );
  Swapper Swapper_171 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_171_io_a0),
    .io_a1(Swapper_171_io_a1),
    .io_z0(Swapper_171_io_z0),
    .io_z1(Swapper_171_io_z1)
  );
  Swapper Swapper_172 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_172_io_a0),
    .io_a1(Swapper_172_io_a1),
    .io_z0(Swapper_172_io_z0),
    .io_z1(Swapper_172_io_z1)
  );
  Swapper Swapper_173 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_173_io_a0),
    .io_a1(Swapper_173_io_a1),
    .io_z0(Swapper_173_io_z0),
    .io_z1(Swapper_173_io_z1)
  );
  Swapper Swapper_174 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_174_io_a0),
    .io_a1(Swapper_174_io_a1),
    .io_z0(Swapper_174_io_z0),
    .io_z1(Swapper_174_io_z1)
  );
  Swapper Swapper_175 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_175_io_a0),
    .io_a1(Swapper_175_io_a1),
    .io_z0(Swapper_175_io_z0),
    .io_z1(Swapper_175_io_z1)
  );
  Swapper Swapper_176 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_176_io_a0),
    .io_a1(Swapper_176_io_a1),
    .io_z0(Swapper_176_io_z0),
    .io_z1(Swapper_176_io_z1)
  );
  Swapper Swapper_177 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_177_io_a0),
    .io_a1(Swapper_177_io_a1),
    .io_z0(Swapper_177_io_z0),
    .io_z1(Swapper_177_io_z1)
  );
  Swapper Swapper_178 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_178_io_a0),
    .io_a1(Swapper_178_io_a1),
    .io_z0(Swapper_178_io_z0),
    .io_z1(Swapper_178_io_z1)
  );
  Swapper Swapper_179 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_179_io_a0),
    .io_a1(Swapper_179_io_a1),
    .io_z0(Swapper_179_io_z0),
    .io_z1(Swapper_179_io_z1)
  );
  Swapper Swapper_180 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_180_io_a0),
    .io_a1(Swapper_180_io_a1),
    .io_z0(Swapper_180_io_z0),
    .io_z1(Swapper_180_io_z1)
  );
  Swapper Swapper_181 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_181_io_a0),
    .io_a1(Swapper_181_io_a1),
    .io_z0(Swapper_181_io_z0),
    .io_z1(Swapper_181_io_z1)
  );
  Swapper Swapper_182 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_182_io_a0),
    .io_a1(Swapper_182_io_a1),
    .io_z0(Swapper_182_io_z0),
    .io_z1(Swapper_182_io_z1)
  );
  Swapper Swapper_183 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_183_io_a0),
    .io_a1(Swapper_183_io_a1),
    .io_z0(Swapper_183_io_z0),
    .io_z1(Swapper_183_io_z1)
  );
  Swapper Swapper_184 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_184_io_a0),
    .io_a1(Swapper_184_io_a1),
    .io_z0(Swapper_184_io_z0),
    .io_z1(Swapper_184_io_z1)
  );
  Swapper Swapper_185 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_185_io_a0),
    .io_a1(Swapper_185_io_a1),
    .io_z0(Swapper_185_io_z0),
    .io_z1(Swapper_185_io_z1)
  );
  Swapper Swapper_186 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_186_io_a0),
    .io_a1(Swapper_186_io_a1),
    .io_z0(Swapper_186_io_z0),
    .io_z1(Swapper_186_io_z1)
  );
  Swapper Swapper_187 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_187_io_a0),
    .io_a1(Swapper_187_io_a1),
    .io_z0(Swapper_187_io_z0),
    .io_z1(Swapper_187_io_z1)
  );
  Swapper Swapper_188 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_188_io_a0),
    .io_a1(Swapper_188_io_a1),
    .io_z0(Swapper_188_io_z0),
    .io_z1(Swapper_188_io_z1)
  );
  Swapper Swapper_189 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_189_io_a0),
    .io_a1(Swapper_189_io_a1),
    .io_z0(Swapper_189_io_z0),
    .io_z1(Swapper_189_io_z1)
  );
  Swapper Swapper_190 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_190_io_a0),
    .io_a1(Swapper_190_io_a1),
    .io_z0(Swapper_190_io_z0),
    .io_z1(Swapper_190_io_z1)
  );
  Swapper Swapper_191 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_191_io_a0),
    .io_a1(Swapper_191_io_a1),
    .io_z0(Swapper_191_io_z0),
    .io_z1(Swapper_191_io_z1)
  );
  Swapper Swapper_192 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_192_io_a0),
    .io_a1(Swapper_192_io_a1),
    .io_z0(Swapper_192_io_z0),
    .io_z1(Swapper_192_io_z1)
  );
  Swapper Swapper_193 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_193_io_a0),
    .io_a1(Swapper_193_io_a1),
    .io_z0(Swapper_193_io_z0),
    .io_z1(Swapper_193_io_z1)
  );
  Swapper Swapper_194 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_194_io_a0),
    .io_a1(Swapper_194_io_a1),
    .io_z0(Swapper_194_io_z0),
    .io_z1(Swapper_194_io_z1)
  );
  Swapper Swapper_195 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_195_io_a0),
    .io_a1(Swapper_195_io_a1),
    .io_z0(Swapper_195_io_z0),
    .io_z1(Swapper_195_io_z1)
  );
  Swapper Swapper_196 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_196_io_a0),
    .io_a1(Swapper_196_io_a1),
    .io_z0(Swapper_196_io_z0),
    .io_z1(Swapper_196_io_z1)
  );
  Swapper Swapper_197 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_197_io_a0),
    .io_a1(Swapper_197_io_a1),
    .io_z0(Swapper_197_io_z0),
    .io_z1(Swapper_197_io_z1)
  );
  Swapper Swapper_198 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_198_io_a0),
    .io_a1(Swapper_198_io_a1),
    .io_z0(Swapper_198_io_z0),
    .io_z1(Swapper_198_io_z1)
  );
  Swapper Swapper_199 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_199_io_a0),
    .io_a1(Swapper_199_io_a1),
    .io_z0(Swapper_199_io_z0),
    .io_z1(Swapper_199_io_z1)
  );
  Swapper Swapper_200 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_200_io_a0),
    .io_a1(Swapper_200_io_a1),
    .io_z0(Swapper_200_io_z0),
    .io_z1(Swapper_200_io_z1)
  );
  Swapper Swapper_201 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_201_io_a0),
    .io_a1(Swapper_201_io_a1),
    .io_z0(Swapper_201_io_z0),
    .io_z1(Swapper_201_io_z1)
  );
  Swapper Swapper_202 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_202_io_a0),
    .io_a1(Swapper_202_io_a1),
    .io_z0(Swapper_202_io_z0),
    .io_z1(Swapper_202_io_z1)
  );
  Swapper Swapper_203 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_203_io_a0),
    .io_a1(Swapper_203_io_a1),
    .io_z0(Swapper_203_io_z0),
    .io_z1(Swapper_203_io_z1)
  );
  Swapper Swapper_204 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_204_io_a0),
    .io_a1(Swapper_204_io_a1),
    .io_z0(Swapper_204_io_z0),
    .io_z1(Swapper_204_io_z1)
  );
  Swapper Swapper_205 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_205_io_a0),
    .io_a1(Swapper_205_io_a1),
    .io_z0(Swapper_205_io_z0),
    .io_z1(Swapper_205_io_z1)
  );
  Swapper Swapper_206 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_206_io_a0),
    .io_a1(Swapper_206_io_a1),
    .io_z0(Swapper_206_io_z0),
    .io_z1(Swapper_206_io_z1)
  );
  Swapper Swapper_207 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_207_io_a0),
    .io_a1(Swapper_207_io_a1),
    .io_z0(Swapper_207_io_z0),
    .io_z1(Swapper_207_io_z1)
  );
  Swapper Swapper_208 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_208_io_a0),
    .io_a1(Swapper_208_io_a1),
    .io_z0(Swapper_208_io_z0),
    .io_z1(Swapper_208_io_z1)
  );
  Swapper Swapper_209 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_209_io_a0),
    .io_a1(Swapper_209_io_a1),
    .io_z0(Swapper_209_io_z0),
    .io_z1(Swapper_209_io_z1)
  );
  Swapper Swapper_210 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_210_io_a0),
    .io_a1(Swapper_210_io_a1),
    .io_z0(Swapper_210_io_z0),
    .io_z1(Swapper_210_io_z1)
  );
  Swapper Swapper_211 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_211_io_a0),
    .io_a1(Swapper_211_io_a1),
    .io_z0(Swapper_211_io_z0),
    .io_z1(Swapper_211_io_z1)
  );
  Swapper Swapper_212 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_212_io_a0),
    .io_a1(Swapper_212_io_a1),
    .io_z0(Swapper_212_io_z0),
    .io_z1(Swapper_212_io_z1)
  );
  Swapper Swapper_213 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_213_io_a0),
    .io_a1(Swapper_213_io_a1),
    .io_z0(Swapper_213_io_z0),
    .io_z1(Swapper_213_io_z1)
  );
  Swapper Swapper_214 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_214_io_a0),
    .io_a1(Swapper_214_io_a1),
    .io_z0(Swapper_214_io_z0),
    .io_z1(Swapper_214_io_z1)
  );
  Swapper Swapper_215 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_215_io_a0),
    .io_a1(Swapper_215_io_a1),
    .io_z0(Swapper_215_io_z0),
    .io_z1(Swapper_215_io_z1)
  );
  Swapper Swapper_216 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_216_io_a0),
    .io_a1(Swapper_216_io_a1),
    .io_z0(Swapper_216_io_z0),
    .io_z1(Swapper_216_io_z1)
  );
  Swapper Swapper_217 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_217_io_a0),
    .io_a1(Swapper_217_io_a1),
    .io_z0(Swapper_217_io_z0),
    .io_z1(Swapper_217_io_z1)
  );
  Swapper Swapper_218 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_218_io_a0),
    .io_a1(Swapper_218_io_a1),
    .io_z0(Swapper_218_io_z0),
    .io_z1(Swapper_218_io_z1)
  );
  Swapper Swapper_219 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_219_io_a0),
    .io_a1(Swapper_219_io_a1),
    .io_z0(Swapper_219_io_z0),
    .io_z1(Swapper_219_io_z1)
  );
  Swapper Swapper_220 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_220_io_a0),
    .io_a1(Swapper_220_io_a1),
    .io_z0(Swapper_220_io_z0),
    .io_z1(Swapper_220_io_z1)
  );
  Swapper Swapper_221 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_221_io_a0),
    .io_a1(Swapper_221_io_a1),
    .io_z0(Swapper_221_io_z0),
    .io_z1(Swapper_221_io_z1)
  );
  Swapper Swapper_222 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_222_io_a0),
    .io_a1(Swapper_222_io_a1),
    .io_z0(Swapper_222_io_z0),
    .io_z1(Swapper_222_io_z1)
  );
  Swapper Swapper_223 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_223_io_a0),
    .io_a1(Swapper_223_io_a1),
    .io_z0(Swapper_223_io_z0),
    .io_z1(Swapper_223_io_z1)
  );
  Swapper Swapper_224 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_224_io_a0),
    .io_a1(Swapper_224_io_a1),
    .io_z0(Swapper_224_io_z0),
    .io_z1(Swapper_224_io_z1)
  );
  Swapper Swapper_225 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_225_io_a0),
    .io_a1(Swapper_225_io_a1),
    .io_z0(Swapper_225_io_z0),
    .io_z1(Swapper_225_io_z1)
  );
  Swapper Swapper_226 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_226_io_a0),
    .io_a1(Swapper_226_io_a1),
    .io_z0(Swapper_226_io_z0),
    .io_z1(Swapper_226_io_z1)
  );
  Swapper Swapper_227 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_227_io_a0),
    .io_a1(Swapper_227_io_a1),
    .io_z0(Swapper_227_io_z0),
    .io_z1(Swapper_227_io_z1)
  );
  Swapper Swapper_228 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_228_io_a0),
    .io_a1(Swapper_228_io_a1),
    .io_z0(Swapper_228_io_z0),
    .io_z1(Swapper_228_io_z1)
  );
  Swapper Swapper_229 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_229_io_a0),
    .io_a1(Swapper_229_io_a1),
    .io_z0(Swapper_229_io_z0),
    .io_z1(Swapper_229_io_z1)
  );
  Swapper Swapper_230 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_230_io_a0),
    .io_a1(Swapper_230_io_a1),
    .io_z0(Swapper_230_io_z0),
    .io_z1(Swapper_230_io_z1)
  );
  Swapper Swapper_231 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_231_io_a0),
    .io_a1(Swapper_231_io_a1),
    .io_z0(Swapper_231_io_z0),
    .io_z1(Swapper_231_io_z1)
  );
  Swapper Swapper_232 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_232_io_a0),
    .io_a1(Swapper_232_io_a1),
    .io_z0(Swapper_232_io_z0),
    .io_z1(Swapper_232_io_z1)
  );
  Swapper Swapper_233 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_233_io_a0),
    .io_a1(Swapper_233_io_a1),
    .io_z0(Swapper_233_io_z0),
    .io_z1(Swapper_233_io_z1)
  );
  Swapper Swapper_234 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_234_io_a0),
    .io_a1(Swapper_234_io_a1),
    .io_z0(Swapper_234_io_z0),
    .io_z1(Swapper_234_io_z1)
  );
  Swapper Swapper_235 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_235_io_a0),
    .io_a1(Swapper_235_io_a1),
    .io_z0(Swapper_235_io_z0),
    .io_z1(Swapper_235_io_z1)
  );
  Swapper Swapper_236 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_236_io_a0),
    .io_a1(Swapper_236_io_a1),
    .io_z0(Swapper_236_io_z0),
    .io_z1(Swapper_236_io_z1)
  );
  Swapper Swapper_237 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_237_io_a0),
    .io_a1(Swapper_237_io_a1),
    .io_z0(Swapper_237_io_z0),
    .io_z1(Swapper_237_io_z1)
  );
  Swapper Swapper_238 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_238_io_a0),
    .io_a1(Swapper_238_io_a1),
    .io_z0(Swapper_238_io_z0),
    .io_z1(Swapper_238_io_z1)
  );
  Swapper Swapper_239 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_239_io_a0),
    .io_a1(Swapper_239_io_a1),
    .io_z0(Swapper_239_io_z0),
    .io_z1(Swapper_239_io_z1)
  );
  Swapper Swapper_240 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_240_io_a0),
    .io_a1(Swapper_240_io_a1),
    .io_z0(Swapper_240_io_z0),
    .io_z1(Swapper_240_io_z1)
  );
  Swapper Swapper_241 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_241_io_a0),
    .io_a1(Swapper_241_io_a1),
    .io_z0(Swapper_241_io_z0),
    .io_z1(Swapper_241_io_z1)
  );
  Swapper Swapper_242 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_242_io_a0),
    .io_a1(Swapper_242_io_a1),
    .io_z0(Swapper_242_io_z0),
    .io_z1(Swapper_242_io_z1)
  );
  Swapper Swapper_243 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_243_io_a0),
    .io_a1(Swapper_243_io_a1),
    .io_z0(Swapper_243_io_z0),
    .io_z1(Swapper_243_io_z1)
  );
  Swapper Swapper_244 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_244_io_a0),
    .io_a1(Swapper_244_io_a1),
    .io_z0(Swapper_244_io_z0),
    .io_z1(Swapper_244_io_z1)
  );
  Swapper Swapper_245 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_245_io_a0),
    .io_a1(Swapper_245_io_a1),
    .io_z0(Swapper_245_io_z0),
    .io_z1(Swapper_245_io_z1)
  );
  Swapper Swapper_246 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_246_io_a0),
    .io_a1(Swapper_246_io_a1),
    .io_z0(Swapper_246_io_z0),
    .io_z1(Swapper_246_io_z1)
  );
  Swapper Swapper_247 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_247_io_a0),
    .io_a1(Swapper_247_io_a1),
    .io_z0(Swapper_247_io_z0),
    .io_z1(Swapper_247_io_z1)
  );
  Swapper Swapper_248 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_248_io_a0),
    .io_a1(Swapper_248_io_a1),
    .io_z0(Swapper_248_io_z0),
    .io_z1(Swapper_248_io_z1)
  );
  Swapper Swapper_249 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_249_io_a0),
    .io_a1(Swapper_249_io_a1),
    .io_z0(Swapper_249_io_z0),
    .io_z1(Swapper_249_io_z1)
  );
  Swapper Swapper_250 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_250_io_a0),
    .io_a1(Swapper_250_io_a1),
    .io_z0(Swapper_250_io_z0),
    .io_z1(Swapper_250_io_z1)
  );
  Swapper Swapper_251 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_251_io_a0),
    .io_a1(Swapper_251_io_a1),
    .io_z0(Swapper_251_io_z0),
    .io_z1(Swapper_251_io_z1)
  );
  Swapper Swapper_252 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_252_io_a0),
    .io_a1(Swapper_252_io_a1),
    .io_z0(Swapper_252_io_z0),
    .io_z1(Swapper_252_io_z1)
  );
  Swapper Swapper_253 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_253_io_a0),
    .io_a1(Swapper_253_io_a1),
    .io_z0(Swapper_253_io_z0),
    .io_z1(Swapper_253_io_z1)
  );
  Swapper Swapper_254 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_254_io_a0),
    .io_a1(Swapper_254_io_a1),
    .io_z0(Swapper_254_io_z0),
    .io_z1(Swapper_254_io_z1)
  );
  Swapper Swapper_255 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_255_io_a0),
    .io_a1(Swapper_255_io_a1),
    .io_z0(Swapper_255_io_z0),
    .io_z1(Swapper_255_io_z1)
  );
  Swapper Swapper_256 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_256_io_a0),
    .io_a1(Swapper_256_io_a1),
    .io_z0(Swapper_256_io_z0),
    .io_z1(Swapper_256_io_z1)
  );
  Swapper Swapper_257 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_257_io_a0),
    .io_a1(Swapper_257_io_a1),
    .io_z0(Swapper_257_io_z0),
    .io_z1(Swapper_257_io_z1)
  );
  Swapper Swapper_258 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_258_io_a0),
    .io_a1(Swapper_258_io_a1),
    .io_z0(Swapper_258_io_z0),
    .io_z1(Swapper_258_io_z1)
  );
  Swapper Swapper_259 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_259_io_a0),
    .io_a1(Swapper_259_io_a1),
    .io_z0(Swapper_259_io_z0),
    .io_z1(Swapper_259_io_z1)
  );
  Swapper Swapper_260 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_260_io_a0),
    .io_a1(Swapper_260_io_a1),
    .io_z0(Swapper_260_io_z0),
    .io_z1(Swapper_260_io_z1)
  );
  Swapper Swapper_261 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_261_io_a0),
    .io_a1(Swapper_261_io_a1),
    .io_z0(Swapper_261_io_z0),
    .io_z1(Swapper_261_io_z1)
  );
  Swapper Swapper_262 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_262_io_a0),
    .io_a1(Swapper_262_io_a1),
    .io_z0(Swapper_262_io_z0),
    .io_z1(Swapper_262_io_z1)
  );
  Swapper Swapper_263 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_263_io_a0),
    .io_a1(Swapper_263_io_a1),
    .io_z0(Swapper_263_io_z0),
    .io_z1(Swapper_263_io_z1)
  );
  Swapper Swapper_264 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_264_io_a0),
    .io_a1(Swapper_264_io_a1),
    .io_z0(Swapper_264_io_z0),
    .io_z1(Swapper_264_io_z1)
  );
  Swapper Swapper_265 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_265_io_a0),
    .io_a1(Swapper_265_io_a1),
    .io_z0(Swapper_265_io_z0),
    .io_z1(Swapper_265_io_z1)
  );
  Swapper Swapper_266 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_266_io_a0),
    .io_a1(Swapper_266_io_a1),
    .io_z0(Swapper_266_io_z0),
    .io_z1(Swapper_266_io_z1)
  );
  Swapper Swapper_267 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_267_io_a0),
    .io_a1(Swapper_267_io_a1),
    .io_z0(Swapper_267_io_z0),
    .io_z1(Swapper_267_io_z1)
  );
  Swapper Swapper_268 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_268_io_a0),
    .io_a1(Swapper_268_io_a1),
    .io_z0(Swapper_268_io_z0),
    .io_z1(Swapper_268_io_z1)
  );
  Swapper Swapper_269 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_269_io_a0),
    .io_a1(Swapper_269_io_a1),
    .io_z0(Swapper_269_io_z0),
    .io_z1(Swapper_269_io_z1)
  );
  Swapper Swapper_270 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_270_io_a0),
    .io_a1(Swapper_270_io_a1),
    .io_z0(Swapper_270_io_z0),
    .io_z1(Swapper_270_io_z1)
  );
  Swapper Swapper_271 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_271_io_a0),
    .io_a1(Swapper_271_io_a1),
    .io_z0(Swapper_271_io_z0),
    .io_z1(Swapper_271_io_z1)
  );
  Swapper Swapper_272 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_272_io_a0),
    .io_a1(Swapper_272_io_a1),
    .io_z0(Swapper_272_io_z0),
    .io_z1(Swapper_272_io_z1)
  );
  Swapper Swapper_273 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_273_io_a0),
    .io_a1(Swapper_273_io_a1),
    .io_z0(Swapper_273_io_z0),
    .io_z1(Swapper_273_io_z1)
  );
  Swapper Swapper_274 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_274_io_a0),
    .io_a1(Swapper_274_io_a1),
    .io_z0(Swapper_274_io_z0),
    .io_z1(Swapper_274_io_z1)
  );
  Swapper Swapper_275 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_275_io_a0),
    .io_a1(Swapper_275_io_a1),
    .io_z0(Swapper_275_io_z0),
    .io_z1(Swapper_275_io_z1)
  );
  Swapper Swapper_276 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_276_io_a0),
    .io_a1(Swapper_276_io_a1),
    .io_z0(Swapper_276_io_z0),
    .io_z1(Swapper_276_io_z1)
  );
  Swapper Swapper_277 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_277_io_a0),
    .io_a1(Swapper_277_io_a1),
    .io_z0(Swapper_277_io_z0),
    .io_z1(Swapper_277_io_z1)
  );
  Swapper Swapper_278 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_278_io_a0),
    .io_a1(Swapper_278_io_a1),
    .io_z0(Swapper_278_io_z0),
    .io_z1(Swapper_278_io_z1)
  );
  Swapper Swapper_279 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_279_io_a0),
    .io_a1(Swapper_279_io_a1),
    .io_z0(Swapper_279_io_z0),
    .io_z1(Swapper_279_io_z1)
  );
  Swapper Swapper_280 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_280_io_a0),
    .io_a1(Swapper_280_io_a1),
    .io_z0(Swapper_280_io_z0),
    .io_z1(Swapper_280_io_z1)
  );
  Swapper Swapper_281 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_281_io_a0),
    .io_a1(Swapper_281_io_a1),
    .io_z0(Swapper_281_io_z0),
    .io_z1(Swapper_281_io_z1)
  );
  Swapper Swapper_282 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_282_io_a0),
    .io_a1(Swapper_282_io_a1),
    .io_z0(Swapper_282_io_z0),
    .io_z1(Swapper_282_io_z1)
  );
  Swapper Swapper_283 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_283_io_a0),
    .io_a1(Swapper_283_io_a1),
    .io_z0(Swapper_283_io_z0),
    .io_z1(Swapper_283_io_z1)
  );
  Swapper Swapper_284 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_284_io_a0),
    .io_a1(Swapper_284_io_a1),
    .io_z0(Swapper_284_io_z0),
    .io_z1(Swapper_284_io_z1)
  );
  Swapper Swapper_285 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_285_io_a0),
    .io_a1(Swapper_285_io_a1),
    .io_z0(Swapper_285_io_z0),
    .io_z1(Swapper_285_io_z1)
  );
  Swapper Swapper_286 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_286_io_a0),
    .io_a1(Swapper_286_io_a1),
    .io_z0(Swapper_286_io_z0),
    .io_z1(Swapper_286_io_z1)
  );
  Swapper Swapper_287 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_287_io_a0),
    .io_a1(Swapper_287_io_a1),
    .io_z0(Swapper_287_io_z0),
    .io_z1(Swapper_287_io_z1)
  );
  Swapper Swapper_288 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_288_io_a0),
    .io_a1(Swapper_288_io_a1),
    .io_z0(Swapper_288_io_z0),
    .io_z1(Swapper_288_io_z1)
  );
  Swapper Swapper_289 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_289_io_a0),
    .io_a1(Swapper_289_io_a1),
    .io_z0(Swapper_289_io_z0),
    .io_z1(Swapper_289_io_z1)
  );
  Swapper Swapper_290 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_290_io_a0),
    .io_a1(Swapper_290_io_a1),
    .io_z0(Swapper_290_io_z0),
    .io_z1(Swapper_290_io_z1)
  );
  Swapper Swapper_291 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_291_io_a0),
    .io_a1(Swapper_291_io_a1),
    .io_z0(Swapper_291_io_z0),
    .io_z1(Swapper_291_io_z1)
  );
  Swapper Swapper_292 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_292_io_a0),
    .io_a1(Swapper_292_io_a1),
    .io_z0(Swapper_292_io_z0),
    .io_z1(Swapper_292_io_z1)
  );
  Swapper Swapper_293 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_293_io_a0),
    .io_a1(Swapper_293_io_a1),
    .io_z0(Swapper_293_io_z0),
    .io_z1(Swapper_293_io_z1)
  );
  Swapper Swapper_294 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_294_io_a0),
    .io_a1(Swapper_294_io_a1),
    .io_z0(Swapper_294_io_z0),
    .io_z1(Swapper_294_io_z1)
  );
  Swapper Swapper_295 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_295_io_a0),
    .io_a1(Swapper_295_io_a1),
    .io_z0(Swapper_295_io_z0),
    .io_z1(Swapper_295_io_z1)
  );
  Swapper Swapper_296 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_296_io_a0),
    .io_a1(Swapper_296_io_a1),
    .io_z0(Swapper_296_io_z0),
    .io_z1(Swapper_296_io_z1)
  );
  Swapper Swapper_297 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_297_io_a0),
    .io_a1(Swapper_297_io_a1),
    .io_z0(Swapper_297_io_z0),
    .io_z1(Swapper_297_io_z1)
  );
  Swapper Swapper_298 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_298_io_a0),
    .io_a1(Swapper_298_io_a1),
    .io_z0(Swapper_298_io_z0),
    .io_z1(Swapper_298_io_z1)
  );
  Swapper Swapper_299 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_299_io_a0),
    .io_a1(Swapper_299_io_a1),
    .io_z0(Swapper_299_io_z0),
    .io_z1(Swapper_299_io_z1)
  );
  Swapper Swapper_300 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_300_io_a0),
    .io_a1(Swapper_300_io_a1),
    .io_z0(Swapper_300_io_z0),
    .io_z1(Swapper_300_io_z1)
  );
  Swapper Swapper_301 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_301_io_a0),
    .io_a1(Swapper_301_io_a1),
    .io_z0(Swapper_301_io_z0),
    .io_z1(Swapper_301_io_z1)
  );
  Swapper Swapper_302 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_302_io_a0),
    .io_a1(Swapper_302_io_a1),
    .io_z0(Swapper_302_io_z0),
    .io_z1(Swapper_302_io_z1)
  );
  Swapper Swapper_303 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_303_io_a0),
    .io_a1(Swapper_303_io_a1),
    .io_z0(Swapper_303_io_z0),
    .io_z1(Swapper_303_io_z1)
  );
  Swapper Swapper_304 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_304_io_a0),
    .io_a1(Swapper_304_io_a1),
    .io_z0(Swapper_304_io_z0),
    .io_z1(Swapper_304_io_z1)
  );
  Swapper Swapper_305 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_305_io_a0),
    .io_a1(Swapper_305_io_a1),
    .io_z0(Swapper_305_io_z0),
    .io_z1(Swapper_305_io_z1)
  );
  Swapper Swapper_306 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_306_io_a0),
    .io_a1(Swapper_306_io_a1),
    .io_z0(Swapper_306_io_z0),
    .io_z1(Swapper_306_io_z1)
  );
  Swapper Swapper_307 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_307_io_a0),
    .io_a1(Swapper_307_io_a1),
    .io_z0(Swapper_307_io_z0),
    .io_z1(Swapper_307_io_z1)
  );
  Swapper Swapper_308 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_308_io_a0),
    .io_a1(Swapper_308_io_a1),
    .io_z0(Swapper_308_io_z0),
    .io_z1(Swapper_308_io_z1)
  );
  Swapper Swapper_309 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_309_io_a0),
    .io_a1(Swapper_309_io_a1),
    .io_z0(Swapper_309_io_z0),
    .io_z1(Swapper_309_io_z1)
  );
  Swapper Swapper_310 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_310_io_a0),
    .io_a1(Swapper_310_io_a1),
    .io_z0(Swapper_310_io_z0),
    .io_z1(Swapper_310_io_z1)
  );
  Swapper Swapper_311 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_311_io_a0),
    .io_a1(Swapper_311_io_a1),
    .io_z0(Swapper_311_io_z0),
    .io_z1(Swapper_311_io_z1)
  );
  Swapper Swapper_312 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_312_io_a0),
    .io_a1(Swapper_312_io_a1),
    .io_z0(Swapper_312_io_z0),
    .io_z1(Swapper_312_io_z1)
  );
  Swapper Swapper_313 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_313_io_a0),
    .io_a1(Swapper_313_io_a1),
    .io_z0(Swapper_313_io_z0),
    .io_z1(Swapper_313_io_z1)
  );
  Swapper Swapper_314 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_314_io_a0),
    .io_a1(Swapper_314_io_a1),
    .io_z0(Swapper_314_io_z0),
    .io_z1(Swapper_314_io_z1)
  );
  Swapper Swapper_315 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_315_io_a0),
    .io_a1(Swapper_315_io_a1),
    .io_z0(Swapper_315_io_z0),
    .io_z1(Swapper_315_io_z1)
  );
  Swapper Swapper_316 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_316_io_a0),
    .io_a1(Swapper_316_io_a1),
    .io_z0(Swapper_316_io_z0),
    .io_z1(Swapper_316_io_z1)
  );
  Swapper Swapper_317 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_317_io_a0),
    .io_a1(Swapper_317_io_a1),
    .io_z0(Swapper_317_io_z0),
    .io_z1(Swapper_317_io_z1)
  );
  Swapper Swapper_318 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_318_io_a0),
    .io_a1(Swapper_318_io_a1),
    .io_z0(Swapper_318_io_z0),
    .io_z1(Swapper_318_io_z1)
  );
  Swapper Swapper_319 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_319_io_a0),
    .io_a1(Swapper_319_io_a1),
    .io_z0(Swapper_319_io_z0),
    .io_z1(Swapper_319_io_z1)
  );
  Swapper Swapper_320 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_320_io_a0),
    .io_a1(Swapper_320_io_a1),
    .io_z0(Swapper_320_io_z0),
    .io_z1(Swapper_320_io_z1)
  );
  Swapper Swapper_321 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_321_io_a0),
    .io_a1(Swapper_321_io_a1),
    .io_z0(Swapper_321_io_z0),
    .io_z1(Swapper_321_io_z1)
  );
  Swapper Swapper_322 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_322_io_a0),
    .io_a1(Swapper_322_io_a1),
    .io_z0(Swapper_322_io_z0),
    .io_z1(Swapper_322_io_z1)
  );
  Swapper Swapper_323 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_323_io_a0),
    .io_a1(Swapper_323_io_a1),
    .io_z0(Swapper_323_io_z0),
    .io_z1(Swapper_323_io_z1)
  );
  Swapper Swapper_324 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_324_io_a0),
    .io_a1(Swapper_324_io_a1),
    .io_z0(Swapper_324_io_z0),
    .io_z1(Swapper_324_io_z1)
  );
  Swapper Swapper_325 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_325_io_a0),
    .io_a1(Swapper_325_io_a1),
    .io_z0(Swapper_325_io_z0),
    .io_z1(Swapper_325_io_z1)
  );
  Swapper Swapper_326 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_326_io_a0),
    .io_a1(Swapper_326_io_a1),
    .io_z0(Swapper_326_io_z0),
    .io_z1(Swapper_326_io_z1)
  );
  Swapper Swapper_327 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_327_io_a0),
    .io_a1(Swapper_327_io_a1),
    .io_z0(Swapper_327_io_z0),
    .io_z1(Swapper_327_io_z1)
  );
  Swapper Swapper_328 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_328_io_a0),
    .io_a1(Swapper_328_io_a1),
    .io_z0(Swapper_328_io_z0),
    .io_z1(Swapper_328_io_z1)
  );
  Swapper Swapper_329 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_329_io_a0),
    .io_a1(Swapper_329_io_a1),
    .io_z0(Swapper_329_io_z0),
    .io_z1(Swapper_329_io_z1)
  );
  Swapper Swapper_330 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_330_io_a0),
    .io_a1(Swapper_330_io_a1),
    .io_z0(Swapper_330_io_z0),
    .io_z1(Swapper_330_io_z1)
  );
  Swapper Swapper_331 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_331_io_a0),
    .io_a1(Swapper_331_io_a1),
    .io_z0(Swapper_331_io_z0),
    .io_z1(Swapper_331_io_z1)
  );
  Swapper Swapper_332 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_332_io_a0),
    .io_a1(Swapper_332_io_a1),
    .io_z0(Swapper_332_io_z0),
    .io_z1(Swapper_332_io_z1)
  );
  Swapper Swapper_333 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_333_io_a0),
    .io_a1(Swapper_333_io_a1),
    .io_z0(Swapper_333_io_z0),
    .io_z1(Swapper_333_io_z1)
  );
  Swapper Swapper_334 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_334_io_a0),
    .io_a1(Swapper_334_io_a1),
    .io_z0(Swapper_334_io_z0),
    .io_z1(Swapper_334_io_z1)
  );
  Swapper Swapper_335 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_335_io_a0),
    .io_a1(Swapper_335_io_a1),
    .io_z0(Swapper_335_io_z0),
    .io_z1(Swapper_335_io_z1)
  );
  Swapper Swapper_336 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_336_io_a0),
    .io_a1(Swapper_336_io_a1),
    .io_z0(Swapper_336_io_z0),
    .io_z1(Swapper_336_io_z1)
  );
  Swapper Swapper_337 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_337_io_a0),
    .io_a1(Swapper_337_io_a1),
    .io_z0(Swapper_337_io_z0),
    .io_z1(Swapper_337_io_z1)
  );
  Swapper Swapper_338 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_338_io_a0),
    .io_a1(Swapper_338_io_a1),
    .io_z0(Swapper_338_io_z0),
    .io_z1(Swapper_338_io_z1)
  );
  Swapper Swapper_339 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_339_io_a0),
    .io_a1(Swapper_339_io_a1),
    .io_z0(Swapper_339_io_z0),
    .io_z1(Swapper_339_io_z1)
  );
  Swapper Swapper_340 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_340_io_a0),
    .io_a1(Swapper_340_io_a1),
    .io_z0(Swapper_340_io_z0),
    .io_z1(Swapper_340_io_z1)
  );
  Swapper Swapper_341 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_341_io_a0),
    .io_a1(Swapper_341_io_a1),
    .io_z0(Swapper_341_io_z0),
    .io_z1(Swapper_341_io_z1)
  );
  Swapper Swapper_342 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_342_io_a0),
    .io_a1(Swapper_342_io_a1),
    .io_z0(Swapper_342_io_z0),
    .io_z1(Swapper_342_io_z1)
  );
  Swapper Swapper_343 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_343_io_a0),
    .io_a1(Swapper_343_io_a1),
    .io_z0(Swapper_343_io_z0),
    .io_z1(Swapper_343_io_z1)
  );
  Swapper Swapper_344 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_344_io_a0),
    .io_a1(Swapper_344_io_a1),
    .io_z0(Swapper_344_io_z0),
    .io_z1(Swapper_344_io_z1)
  );
  Swapper Swapper_345 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_345_io_a0),
    .io_a1(Swapper_345_io_a1),
    .io_z0(Swapper_345_io_z0),
    .io_z1(Swapper_345_io_z1)
  );
  Swapper Swapper_346 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_346_io_a0),
    .io_a1(Swapper_346_io_a1),
    .io_z0(Swapper_346_io_z0),
    .io_z1(Swapper_346_io_z1)
  );
  Swapper Swapper_347 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_347_io_a0),
    .io_a1(Swapper_347_io_a1),
    .io_z0(Swapper_347_io_z0),
    .io_z1(Swapper_347_io_z1)
  );
  Swapper Swapper_348 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_348_io_a0),
    .io_a1(Swapper_348_io_a1),
    .io_z0(Swapper_348_io_z0),
    .io_z1(Swapper_348_io_z1)
  );
  Swapper Swapper_349 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_349_io_a0),
    .io_a1(Swapper_349_io_a1),
    .io_z0(Swapper_349_io_z0),
    .io_z1(Swapper_349_io_z1)
  );
  Swapper Swapper_350 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_350_io_a0),
    .io_a1(Swapper_350_io_a1),
    .io_z0(Swapper_350_io_z0),
    .io_z1(Swapper_350_io_z1)
  );
  Swapper Swapper_351 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_351_io_a0),
    .io_a1(Swapper_351_io_a1),
    .io_z0(Swapper_351_io_z0),
    .io_z1(Swapper_351_io_z1)
  );
  Swapper Swapper_352 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_352_io_a0),
    .io_a1(Swapper_352_io_a1),
    .io_z0(Swapper_352_io_z0),
    .io_z1(Swapper_352_io_z1)
  );
  Swapper Swapper_353 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_353_io_a0),
    .io_a1(Swapper_353_io_a1),
    .io_z0(Swapper_353_io_z0),
    .io_z1(Swapper_353_io_z1)
  );
  Swapper Swapper_354 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_354_io_a0),
    .io_a1(Swapper_354_io_a1),
    .io_z0(Swapper_354_io_z0),
    .io_z1(Swapper_354_io_z1)
  );
  Swapper Swapper_355 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_355_io_a0),
    .io_a1(Swapper_355_io_a1),
    .io_z0(Swapper_355_io_z0),
    .io_z1(Swapper_355_io_z1)
  );
  Swapper Swapper_356 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_356_io_a0),
    .io_a1(Swapper_356_io_a1),
    .io_z0(Swapper_356_io_z0),
    .io_z1(Swapper_356_io_z1)
  );
  Swapper Swapper_357 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_357_io_a0),
    .io_a1(Swapper_357_io_a1),
    .io_z0(Swapper_357_io_z0),
    .io_z1(Swapper_357_io_z1)
  );
  Swapper Swapper_358 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_358_io_a0),
    .io_a1(Swapper_358_io_a1),
    .io_z0(Swapper_358_io_z0),
    .io_z1(Swapper_358_io_z1)
  );
  Swapper Swapper_359 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_359_io_a0),
    .io_a1(Swapper_359_io_a1),
    .io_z0(Swapper_359_io_z0),
    .io_z1(Swapper_359_io_z1)
  );
  Swapper Swapper_360 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_360_io_a0),
    .io_a1(Swapper_360_io_a1),
    .io_z0(Swapper_360_io_z0),
    .io_z1(Swapper_360_io_z1)
  );
  Swapper Swapper_361 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_361_io_a0),
    .io_a1(Swapper_361_io_a1),
    .io_z0(Swapper_361_io_z0),
    .io_z1(Swapper_361_io_z1)
  );
  Swapper Swapper_362 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_362_io_a0),
    .io_a1(Swapper_362_io_a1),
    .io_z0(Swapper_362_io_z0),
    .io_z1(Swapper_362_io_z1)
  );
  Swapper Swapper_363 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_363_io_a0),
    .io_a1(Swapper_363_io_a1),
    .io_z0(Swapper_363_io_z0),
    .io_z1(Swapper_363_io_z1)
  );
  Swapper Swapper_364 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_364_io_a0),
    .io_a1(Swapper_364_io_a1),
    .io_z0(Swapper_364_io_z0),
    .io_z1(Swapper_364_io_z1)
  );
  Swapper Swapper_365 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_365_io_a0),
    .io_a1(Swapper_365_io_a1),
    .io_z0(Swapper_365_io_z0),
    .io_z1(Swapper_365_io_z1)
  );
  Swapper Swapper_366 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_366_io_a0),
    .io_a1(Swapper_366_io_a1),
    .io_z0(Swapper_366_io_z0),
    .io_z1(Swapper_366_io_z1)
  );
  Swapper Swapper_367 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_367_io_a0),
    .io_a1(Swapper_367_io_a1),
    .io_z0(Swapper_367_io_z0),
    .io_z1(Swapper_367_io_z1)
  );
  Swapper Swapper_368 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_368_io_a0),
    .io_a1(Swapper_368_io_a1),
    .io_z0(Swapper_368_io_z0),
    .io_z1(Swapper_368_io_z1)
  );
  Swapper Swapper_369 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_369_io_a0),
    .io_a1(Swapper_369_io_a1),
    .io_z0(Swapper_369_io_z0),
    .io_z1(Swapper_369_io_z1)
  );
  Swapper Swapper_370 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_370_io_a0),
    .io_a1(Swapper_370_io_a1),
    .io_z0(Swapper_370_io_z0),
    .io_z1(Swapper_370_io_z1)
  );
  Swapper Swapper_371 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_371_io_a0),
    .io_a1(Swapper_371_io_a1),
    .io_z0(Swapper_371_io_z0),
    .io_z1(Swapper_371_io_z1)
  );
  Swapper Swapper_372 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_372_io_a0),
    .io_a1(Swapper_372_io_a1),
    .io_z0(Swapper_372_io_z0),
    .io_z1(Swapper_372_io_z1)
  );
  Swapper Swapper_373 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_373_io_a0),
    .io_a1(Swapper_373_io_a1),
    .io_z0(Swapper_373_io_z0),
    .io_z1(Swapper_373_io_z1)
  );
  Swapper Swapper_374 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_374_io_a0),
    .io_a1(Swapper_374_io_a1),
    .io_z0(Swapper_374_io_z0),
    .io_z1(Swapper_374_io_z1)
  );
  Swapper Swapper_375 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_375_io_a0),
    .io_a1(Swapper_375_io_a1),
    .io_z0(Swapper_375_io_z0),
    .io_z1(Swapper_375_io_z1)
  );
  Swapper Swapper_376 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_376_io_a0),
    .io_a1(Swapper_376_io_a1),
    .io_z0(Swapper_376_io_z0),
    .io_z1(Swapper_376_io_z1)
  );
  Swapper Swapper_377 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_377_io_a0),
    .io_a1(Swapper_377_io_a1),
    .io_z0(Swapper_377_io_z0),
    .io_z1(Swapper_377_io_z1)
  );
  Swapper Swapper_378 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_378_io_a0),
    .io_a1(Swapper_378_io_a1),
    .io_z0(Swapper_378_io_z0),
    .io_z1(Swapper_378_io_z1)
  );
  Swapper Swapper_379 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_379_io_a0),
    .io_a1(Swapper_379_io_a1),
    .io_z0(Swapper_379_io_z0),
    .io_z1(Swapper_379_io_z1)
  );
  Swapper Swapper_380 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_380_io_a0),
    .io_a1(Swapper_380_io_a1),
    .io_z0(Swapper_380_io_z0),
    .io_z1(Swapper_380_io_z1)
  );
  Swapper Swapper_381 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_381_io_a0),
    .io_a1(Swapper_381_io_a1),
    .io_z0(Swapper_381_io_z0),
    .io_z1(Swapper_381_io_z1)
  );
  Swapper Swapper_382 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_382_io_a0),
    .io_a1(Swapper_382_io_a1),
    .io_z0(Swapper_382_io_z0),
    .io_z1(Swapper_382_io_z1)
  );
  Swapper Swapper_383 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_383_io_a0),
    .io_a1(Swapper_383_io_a1),
    .io_z0(Swapper_383_io_z0),
    .io_z1(Swapper_383_io_z1)
  );
  Swapper Swapper_384 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_384_io_a0),
    .io_a1(Swapper_384_io_a1),
    .io_z0(Swapper_384_io_z0),
    .io_z1(Swapper_384_io_z1)
  );
  Swapper Swapper_385 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_385_io_a0),
    .io_a1(Swapper_385_io_a1),
    .io_z0(Swapper_385_io_z0),
    .io_z1(Swapper_385_io_z1)
  );
  Swapper Swapper_386 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_386_io_a0),
    .io_a1(Swapper_386_io_a1),
    .io_z0(Swapper_386_io_z0),
    .io_z1(Swapper_386_io_z1)
  );
  Swapper Swapper_387 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_387_io_a0),
    .io_a1(Swapper_387_io_a1),
    .io_z0(Swapper_387_io_z0),
    .io_z1(Swapper_387_io_z1)
  );
  Swapper Swapper_388 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_388_io_a0),
    .io_a1(Swapper_388_io_a1),
    .io_z0(Swapper_388_io_z0),
    .io_z1(Swapper_388_io_z1)
  );
  Swapper Swapper_389 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_389_io_a0),
    .io_a1(Swapper_389_io_a1),
    .io_z0(Swapper_389_io_z0),
    .io_z1(Swapper_389_io_z1)
  );
  Swapper Swapper_390 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_390_io_a0),
    .io_a1(Swapper_390_io_a1),
    .io_z0(Swapper_390_io_z0),
    .io_z1(Swapper_390_io_z1)
  );
  Swapper Swapper_391 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_391_io_a0),
    .io_a1(Swapper_391_io_a1),
    .io_z0(Swapper_391_io_z0),
    .io_z1(Swapper_391_io_z1)
  );
  Swapper Swapper_392 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_392_io_a0),
    .io_a1(Swapper_392_io_a1),
    .io_z0(Swapper_392_io_z0),
    .io_z1(Swapper_392_io_z1)
  );
  Swapper Swapper_393 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_393_io_a0),
    .io_a1(Swapper_393_io_a1),
    .io_z0(Swapper_393_io_z0),
    .io_z1(Swapper_393_io_z1)
  );
  Swapper Swapper_394 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_394_io_a0),
    .io_a1(Swapper_394_io_a1),
    .io_z0(Swapper_394_io_z0),
    .io_z1(Swapper_394_io_z1)
  );
  Swapper Swapper_395 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_395_io_a0),
    .io_a1(Swapper_395_io_a1),
    .io_z0(Swapper_395_io_z0),
    .io_z1(Swapper_395_io_z1)
  );
  Swapper Swapper_396 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_396_io_a0),
    .io_a1(Swapper_396_io_a1),
    .io_z0(Swapper_396_io_z0),
    .io_z1(Swapper_396_io_z1)
  );
  Swapper Swapper_397 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_397_io_a0),
    .io_a1(Swapper_397_io_a1),
    .io_z0(Swapper_397_io_z0),
    .io_z1(Swapper_397_io_z1)
  );
  Swapper Swapper_398 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_398_io_a0),
    .io_a1(Swapper_398_io_a1),
    .io_z0(Swapper_398_io_z0),
    .io_z1(Swapper_398_io_z1)
  );
  Swapper Swapper_399 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_399_io_a0),
    .io_a1(Swapper_399_io_a1),
    .io_z0(Swapper_399_io_z0),
    .io_z1(Swapper_399_io_z1)
  );
  Swapper Swapper_400 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_400_io_a0),
    .io_a1(Swapper_400_io_a1),
    .io_z0(Swapper_400_io_z0),
    .io_z1(Swapper_400_io_z1)
  );
  Swapper Swapper_401 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_401_io_a0),
    .io_a1(Swapper_401_io_a1),
    .io_z0(Swapper_401_io_z0),
    .io_z1(Swapper_401_io_z1)
  );
  Swapper Swapper_402 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_402_io_a0),
    .io_a1(Swapper_402_io_a1),
    .io_z0(Swapper_402_io_z0),
    .io_z1(Swapper_402_io_z1)
  );
  Swapper Swapper_403 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_403_io_a0),
    .io_a1(Swapper_403_io_a1),
    .io_z0(Swapper_403_io_z0),
    .io_z1(Swapper_403_io_z1)
  );
  Swapper Swapper_404 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_404_io_a0),
    .io_a1(Swapper_404_io_a1),
    .io_z0(Swapper_404_io_z0),
    .io_z1(Swapper_404_io_z1)
  );
  Swapper Swapper_405 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_405_io_a0),
    .io_a1(Swapper_405_io_a1),
    .io_z0(Swapper_405_io_z0),
    .io_z1(Swapper_405_io_z1)
  );
  Swapper Swapper_406 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_406_io_a0),
    .io_a1(Swapper_406_io_a1),
    .io_z0(Swapper_406_io_z0),
    .io_z1(Swapper_406_io_z1)
  );
  Swapper Swapper_407 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_407_io_a0),
    .io_a1(Swapper_407_io_a1),
    .io_z0(Swapper_407_io_z0),
    .io_z1(Swapper_407_io_z1)
  );
  Swapper Swapper_408 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_408_io_a0),
    .io_a1(Swapper_408_io_a1),
    .io_z0(Swapper_408_io_z0),
    .io_z1(Swapper_408_io_z1)
  );
  Swapper Swapper_409 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_409_io_a0),
    .io_a1(Swapper_409_io_a1),
    .io_z0(Swapper_409_io_z0),
    .io_z1(Swapper_409_io_z1)
  );
  Swapper Swapper_410 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_410_io_a0),
    .io_a1(Swapper_410_io_a1),
    .io_z0(Swapper_410_io_z0),
    .io_z1(Swapper_410_io_z1)
  );
  Swapper Swapper_411 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_411_io_a0),
    .io_a1(Swapper_411_io_a1),
    .io_z0(Swapper_411_io_z0),
    .io_z1(Swapper_411_io_z1)
  );
  Swapper Swapper_412 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_412_io_a0),
    .io_a1(Swapper_412_io_a1),
    .io_z0(Swapper_412_io_z0),
    .io_z1(Swapper_412_io_z1)
  );
  Swapper Swapper_413 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_413_io_a0),
    .io_a1(Swapper_413_io_a1),
    .io_z0(Swapper_413_io_z0),
    .io_z1(Swapper_413_io_z1)
  );
  Swapper Swapper_414 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_414_io_a0),
    .io_a1(Swapper_414_io_a1),
    .io_z0(Swapper_414_io_z0),
    .io_z1(Swapper_414_io_z1)
  );
  Swapper Swapper_415 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_415_io_a0),
    .io_a1(Swapper_415_io_a1),
    .io_z0(Swapper_415_io_z0),
    .io_z1(Swapper_415_io_z1)
  );
  Swapper Swapper_416 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_416_io_a0),
    .io_a1(Swapper_416_io_a1),
    .io_z0(Swapper_416_io_z0),
    .io_z1(Swapper_416_io_z1)
  );
  Swapper Swapper_417 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_417_io_a0),
    .io_a1(Swapper_417_io_a1),
    .io_z0(Swapper_417_io_z0),
    .io_z1(Swapper_417_io_z1)
  );
  Swapper Swapper_418 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_418_io_a0),
    .io_a1(Swapper_418_io_a1),
    .io_z0(Swapper_418_io_z0),
    .io_z1(Swapper_418_io_z1)
  );
  Swapper Swapper_419 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_419_io_a0),
    .io_a1(Swapper_419_io_a1),
    .io_z0(Swapper_419_io_z0),
    .io_z1(Swapper_419_io_z1)
  );
  Swapper Swapper_420 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_420_io_a0),
    .io_a1(Swapper_420_io_a1),
    .io_z0(Swapper_420_io_z0),
    .io_z1(Swapper_420_io_z1)
  );
  Swapper Swapper_421 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_421_io_a0),
    .io_a1(Swapper_421_io_a1),
    .io_z0(Swapper_421_io_z0),
    .io_z1(Swapper_421_io_z1)
  );
  Swapper Swapper_422 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_422_io_a0),
    .io_a1(Swapper_422_io_a1),
    .io_z0(Swapper_422_io_z0),
    .io_z1(Swapper_422_io_z1)
  );
  Swapper Swapper_423 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_423_io_a0),
    .io_a1(Swapper_423_io_a1),
    .io_z0(Swapper_423_io_z0),
    .io_z1(Swapper_423_io_z1)
  );
  Swapper Swapper_424 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_424_io_a0),
    .io_a1(Swapper_424_io_a1),
    .io_z0(Swapper_424_io_z0),
    .io_z1(Swapper_424_io_z1)
  );
  Swapper Swapper_425 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_425_io_a0),
    .io_a1(Swapper_425_io_a1),
    .io_z0(Swapper_425_io_z0),
    .io_z1(Swapper_425_io_z1)
  );
  Swapper Swapper_426 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_426_io_a0),
    .io_a1(Swapper_426_io_a1),
    .io_z0(Swapper_426_io_z0),
    .io_z1(Swapper_426_io_z1)
  );
  Swapper Swapper_427 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_427_io_a0),
    .io_a1(Swapper_427_io_a1),
    .io_z0(Swapper_427_io_z0),
    .io_z1(Swapper_427_io_z1)
  );
  Swapper Swapper_428 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_428_io_a0),
    .io_a1(Swapper_428_io_a1),
    .io_z0(Swapper_428_io_z0),
    .io_z1(Swapper_428_io_z1)
  );
  Swapper Swapper_429 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_429_io_a0),
    .io_a1(Swapper_429_io_a1),
    .io_z0(Swapper_429_io_z0),
    .io_z1(Swapper_429_io_z1)
  );
  Swapper Swapper_430 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_430_io_a0),
    .io_a1(Swapper_430_io_a1),
    .io_z0(Swapper_430_io_z0),
    .io_z1(Swapper_430_io_z1)
  );
  Swapper Swapper_431 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_431_io_a0),
    .io_a1(Swapper_431_io_a1),
    .io_z0(Swapper_431_io_z0),
    .io_z1(Swapper_431_io_z1)
  );
  Swapper Swapper_432 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_432_io_a0),
    .io_a1(Swapper_432_io_a1),
    .io_z0(Swapper_432_io_z0),
    .io_z1(Swapper_432_io_z1)
  );
  Swapper Swapper_433 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_433_io_a0),
    .io_a1(Swapper_433_io_a1),
    .io_z0(Swapper_433_io_z0),
    .io_z1(Swapper_433_io_z1)
  );
  Swapper Swapper_434 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_434_io_a0),
    .io_a1(Swapper_434_io_a1),
    .io_z0(Swapper_434_io_z0),
    .io_z1(Swapper_434_io_z1)
  );
  Swapper Swapper_435 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_435_io_a0),
    .io_a1(Swapper_435_io_a1),
    .io_z0(Swapper_435_io_z0),
    .io_z1(Swapper_435_io_z1)
  );
  Swapper Swapper_436 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_436_io_a0),
    .io_a1(Swapper_436_io_a1),
    .io_z0(Swapper_436_io_z0),
    .io_z1(Swapper_436_io_z1)
  );
  Swapper Swapper_437 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_437_io_a0),
    .io_a1(Swapper_437_io_a1),
    .io_z0(Swapper_437_io_z0),
    .io_z1(Swapper_437_io_z1)
  );
  Swapper Swapper_438 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_438_io_a0),
    .io_a1(Swapper_438_io_a1),
    .io_z0(Swapper_438_io_z0),
    .io_z1(Swapper_438_io_z1)
  );
  Swapper Swapper_439 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_439_io_a0),
    .io_a1(Swapper_439_io_a1),
    .io_z0(Swapper_439_io_z0),
    .io_z1(Swapper_439_io_z1)
  );
  Swapper Swapper_440 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_440_io_a0),
    .io_a1(Swapper_440_io_a1),
    .io_z0(Swapper_440_io_z0),
    .io_z1(Swapper_440_io_z1)
  );
  Swapper Swapper_441 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_441_io_a0),
    .io_a1(Swapper_441_io_a1),
    .io_z0(Swapper_441_io_z0),
    .io_z1(Swapper_441_io_z1)
  );
  Swapper Swapper_442 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_442_io_a0),
    .io_a1(Swapper_442_io_a1),
    .io_z0(Swapper_442_io_z0),
    .io_z1(Swapper_442_io_z1)
  );
  Swapper Swapper_443 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_443_io_a0),
    .io_a1(Swapper_443_io_a1),
    .io_z0(Swapper_443_io_z0),
    .io_z1(Swapper_443_io_z1)
  );
  Swapper Swapper_444 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_444_io_a0),
    .io_a1(Swapper_444_io_a1),
    .io_z0(Swapper_444_io_z0),
    .io_z1(Swapper_444_io_z1)
  );
  Swapper Swapper_445 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_445_io_a0),
    .io_a1(Swapper_445_io_a1),
    .io_z0(Swapper_445_io_z0),
    .io_z1(Swapper_445_io_z1)
  );
  Swapper Swapper_446 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_446_io_a0),
    .io_a1(Swapper_446_io_a1),
    .io_z0(Swapper_446_io_z0),
    .io_z1(Swapper_446_io_z1)
  );
  Swapper Swapper_447 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_447_io_a0),
    .io_a1(Swapper_447_io_a1),
    .io_z0(Swapper_447_io_z0),
    .io_z1(Swapper_447_io_z1)
  );
  Swapper Swapper_448 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_448_io_a0),
    .io_a1(Swapper_448_io_a1),
    .io_z0(Swapper_448_io_z0),
    .io_z1(Swapper_448_io_z1)
  );
  Swapper Swapper_449 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_449_io_a0),
    .io_a1(Swapper_449_io_a1),
    .io_z0(Swapper_449_io_z0),
    .io_z1(Swapper_449_io_z1)
  );
  Swapper Swapper_450 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_450_io_a0),
    .io_a1(Swapper_450_io_a1),
    .io_z0(Swapper_450_io_z0),
    .io_z1(Swapper_450_io_z1)
  );
  Swapper Swapper_451 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_451_io_a0),
    .io_a1(Swapper_451_io_a1),
    .io_z0(Swapper_451_io_z0),
    .io_z1(Swapper_451_io_z1)
  );
  Swapper Swapper_452 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_452_io_a0),
    .io_a1(Swapper_452_io_a1),
    .io_z0(Swapper_452_io_z0),
    .io_z1(Swapper_452_io_z1)
  );
  Swapper Swapper_453 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_453_io_a0),
    .io_a1(Swapper_453_io_a1),
    .io_z0(Swapper_453_io_z0),
    .io_z1(Swapper_453_io_z1)
  );
  Swapper Swapper_454 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_454_io_a0),
    .io_a1(Swapper_454_io_a1),
    .io_z0(Swapper_454_io_z0),
    .io_z1(Swapper_454_io_z1)
  );
  Swapper Swapper_455 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_455_io_a0),
    .io_a1(Swapper_455_io_a1),
    .io_z0(Swapper_455_io_z0),
    .io_z1(Swapper_455_io_z1)
  );
  Swapper Swapper_456 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_456_io_a0),
    .io_a1(Swapper_456_io_a1),
    .io_z0(Swapper_456_io_z0),
    .io_z1(Swapper_456_io_z1)
  );
  Swapper Swapper_457 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_457_io_a0),
    .io_a1(Swapper_457_io_a1),
    .io_z0(Swapper_457_io_z0),
    .io_z1(Swapper_457_io_z1)
  );
  Swapper Swapper_458 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_458_io_a0),
    .io_a1(Swapper_458_io_a1),
    .io_z0(Swapper_458_io_z0),
    .io_z1(Swapper_458_io_z1)
  );
  Swapper Swapper_459 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_459_io_a0),
    .io_a1(Swapper_459_io_a1),
    .io_z0(Swapper_459_io_z0),
    .io_z1(Swapper_459_io_z1)
  );
  Swapper Swapper_460 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_460_io_a0),
    .io_a1(Swapper_460_io_a1),
    .io_z0(Swapper_460_io_z0),
    .io_z1(Swapper_460_io_z1)
  );
  Swapper Swapper_461 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_461_io_a0),
    .io_a1(Swapper_461_io_a1),
    .io_z0(Swapper_461_io_z0),
    .io_z1(Swapper_461_io_z1)
  );
  Swapper Swapper_462 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_462_io_a0),
    .io_a1(Swapper_462_io_a1),
    .io_z0(Swapper_462_io_z0),
    .io_z1(Swapper_462_io_z1)
  );
  Swapper Swapper_463 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_463_io_a0),
    .io_a1(Swapper_463_io_a1),
    .io_z0(Swapper_463_io_z0),
    .io_z1(Swapper_463_io_z1)
  );
  Swapper Swapper_464 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_464_io_a0),
    .io_a1(Swapper_464_io_a1),
    .io_z0(Swapper_464_io_z0),
    .io_z1(Swapper_464_io_z1)
  );
  Swapper Swapper_465 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_465_io_a0),
    .io_a1(Swapper_465_io_a1),
    .io_z0(Swapper_465_io_z0),
    .io_z1(Swapper_465_io_z1)
  );
  Swapper Swapper_466 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_466_io_a0),
    .io_a1(Swapper_466_io_a1),
    .io_z0(Swapper_466_io_z0),
    .io_z1(Swapper_466_io_z1)
  );
  Swapper Swapper_467 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_467_io_a0),
    .io_a1(Swapper_467_io_a1),
    .io_z0(Swapper_467_io_z0),
    .io_z1(Swapper_467_io_z1)
  );
  Swapper Swapper_468 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_468_io_a0),
    .io_a1(Swapper_468_io_a1),
    .io_z0(Swapper_468_io_z0),
    .io_z1(Swapper_468_io_z1)
  );
  Swapper Swapper_469 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_469_io_a0),
    .io_a1(Swapper_469_io_a1),
    .io_z0(Swapper_469_io_z0),
    .io_z1(Swapper_469_io_z1)
  );
  Swapper Swapper_470 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_470_io_a0),
    .io_a1(Swapper_470_io_a1),
    .io_z0(Swapper_470_io_z0),
    .io_z1(Swapper_470_io_z1)
  );
  Swapper Swapper_471 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_471_io_a0),
    .io_a1(Swapper_471_io_a1),
    .io_z0(Swapper_471_io_z0),
    .io_z1(Swapper_471_io_z1)
  );
  Swapper Swapper_472 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_472_io_a0),
    .io_a1(Swapper_472_io_a1),
    .io_z0(Swapper_472_io_z0),
    .io_z1(Swapper_472_io_z1)
  );
  Swapper Swapper_473 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_473_io_a0),
    .io_a1(Swapper_473_io_a1),
    .io_z0(Swapper_473_io_z0),
    .io_z1(Swapper_473_io_z1)
  );
  Swapper Swapper_474 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_474_io_a0),
    .io_a1(Swapper_474_io_a1),
    .io_z0(Swapper_474_io_z0),
    .io_z1(Swapper_474_io_z1)
  );
  Swapper Swapper_475 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_475_io_a0),
    .io_a1(Swapper_475_io_a1),
    .io_z0(Swapper_475_io_z0),
    .io_z1(Swapper_475_io_z1)
  );
  Swapper Swapper_476 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_476_io_a0),
    .io_a1(Swapper_476_io_a1),
    .io_z0(Swapper_476_io_z0),
    .io_z1(Swapper_476_io_z1)
  );
  Swapper Swapper_477 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_477_io_a0),
    .io_a1(Swapper_477_io_a1),
    .io_z0(Swapper_477_io_z0),
    .io_z1(Swapper_477_io_z1)
  );
  Swapper Swapper_478 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_478_io_a0),
    .io_a1(Swapper_478_io_a1),
    .io_z0(Swapper_478_io_z0),
    .io_z1(Swapper_478_io_z1)
  );
  Swapper Swapper_479 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_479_io_a0),
    .io_a1(Swapper_479_io_a1),
    .io_z0(Swapper_479_io_z0),
    .io_z1(Swapper_479_io_z1)
  );
  Swapper Swapper_480 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_480_io_a0),
    .io_a1(Swapper_480_io_a1),
    .io_z0(Swapper_480_io_z0),
    .io_z1(Swapper_480_io_z1)
  );
  Swapper Swapper_481 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_481_io_a0),
    .io_a1(Swapper_481_io_a1),
    .io_z0(Swapper_481_io_z0),
    .io_z1(Swapper_481_io_z1)
  );
  Swapper Swapper_482 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_482_io_a0),
    .io_a1(Swapper_482_io_a1),
    .io_z0(Swapper_482_io_z0),
    .io_z1(Swapper_482_io_z1)
  );
  Swapper Swapper_483 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_483_io_a0),
    .io_a1(Swapper_483_io_a1),
    .io_z0(Swapper_483_io_z0),
    .io_z1(Swapper_483_io_z1)
  );
  Swapper Swapper_484 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_484_io_a0),
    .io_a1(Swapper_484_io_a1),
    .io_z0(Swapper_484_io_z0),
    .io_z1(Swapper_484_io_z1)
  );
  Swapper Swapper_485 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_485_io_a0),
    .io_a1(Swapper_485_io_a1),
    .io_z0(Swapper_485_io_z0),
    .io_z1(Swapper_485_io_z1)
  );
  Swapper Swapper_486 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_486_io_a0),
    .io_a1(Swapper_486_io_a1),
    .io_z0(Swapper_486_io_z0),
    .io_z1(Swapper_486_io_z1)
  );
  Swapper Swapper_487 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_487_io_a0),
    .io_a1(Swapper_487_io_a1),
    .io_z0(Swapper_487_io_z0),
    .io_z1(Swapper_487_io_z1)
  );
  Swapper Swapper_488 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_488_io_a0),
    .io_a1(Swapper_488_io_a1),
    .io_z0(Swapper_488_io_z0),
    .io_z1(Swapper_488_io_z1)
  );
  Swapper Swapper_489 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_489_io_a0),
    .io_a1(Swapper_489_io_a1),
    .io_z0(Swapper_489_io_z0),
    .io_z1(Swapper_489_io_z1)
  );
  Swapper Swapper_490 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_490_io_a0),
    .io_a1(Swapper_490_io_a1),
    .io_z0(Swapper_490_io_z0),
    .io_z1(Swapper_490_io_z1)
  );
  Swapper Swapper_491 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_491_io_a0),
    .io_a1(Swapper_491_io_a1),
    .io_z0(Swapper_491_io_z0),
    .io_z1(Swapper_491_io_z1)
  );
  Swapper Swapper_492 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_492_io_a0),
    .io_a1(Swapper_492_io_a1),
    .io_z0(Swapper_492_io_z0),
    .io_z1(Swapper_492_io_z1)
  );
  Swapper Swapper_493 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_493_io_a0),
    .io_a1(Swapper_493_io_a1),
    .io_z0(Swapper_493_io_z0),
    .io_z1(Swapper_493_io_z1)
  );
  Swapper Swapper_494 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_494_io_a0),
    .io_a1(Swapper_494_io_a1),
    .io_z0(Swapper_494_io_z0),
    .io_z1(Swapper_494_io_z1)
  );
  Swapper Swapper_495 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_495_io_a0),
    .io_a1(Swapper_495_io_a1),
    .io_z0(Swapper_495_io_z0),
    .io_z1(Swapper_495_io_z1)
  );
  Swapper Swapper_496 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_496_io_a0),
    .io_a1(Swapper_496_io_a1),
    .io_z0(Swapper_496_io_z0),
    .io_z1(Swapper_496_io_z1)
  );
  Swapper Swapper_497 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_497_io_a0),
    .io_a1(Swapper_497_io_a1),
    .io_z0(Swapper_497_io_z0),
    .io_z1(Swapper_497_io_z1)
  );
  Swapper Swapper_498 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_498_io_a0),
    .io_a1(Swapper_498_io_a1),
    .io_z0(Swapper_498_io_z0),
    .io_z1(Swapper_498_io_z1)
  );
  Swapper Swapper_499 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_499_io_a0),
    .io_a1(Swapper_499_io_a1),
    .io_z0(Swapper_499_io_z0),
    .io_z1(Swapper_499_io_z1)
  );
  Swapper Swapper_500 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_500_io_a0),
    .io_a1(Swapper_500_io_a1),
    .io_z0(Swapper_500_io_z0),
    .io_z1(Swapper_500_io_z1)
  );
  Swapper Swapper_501 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_501_io_a0),
    .io_a1(Swapper_501_io_a1),
    .io_z0(Swapper_501_io_z0),
    .io_z1(Swapper_501_io_z1)
  );
  Swapper Swapper_502 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_502_io_a0),
    .io_a1(Swapper_502_io_a1),
    .io_z0(Swapper_502_io_z0),
    .io_z1(Swapper_502_io_z1)
  );
  Swapper Swapper_503 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_503_io_a0),
    .io_a1(Swapper_503_io_a1),
    .io_z0(Swapper_503_io_z0),
    .io_z1(Swapper_503_io_z1)
  );
  Swapper Swapper_504 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_504_io_a0),
    .io_a1(Swapper_504_io_a1),
    .io_z0(Swapper_504_io_z0),
    .io_z1(Swapper_504_io_z1)
  );
  Swapper Swapper_505 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_505_io_a0),
    .io_a1(Swapper_505_io_a1),
    .io_z0(Swapper_505_io_z0),
    .io_z1(Swapper_505_io_z1)
  );
  Swapper Swapper_506 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_506_io_a0),
    .io_a1(Swapper_506_io_a1),
    .io_z0(Swapper_506_io_z0),
    .io_z1(Swapper_506_io_z1)
  );
  Swapper Swapper_507 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_507_io_a0),
    .io_a1(Swapper_507_io_a1),
    .io_z0(Swapper_507_io_z0),
    .io_z1(Swapper_507_io_z1)
  );
  Swapper Swapper_508 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_508_io_a0),
    .io_a1(Swapper_508_io_a1),
    .io_z0(Swapper_508_io_z0),
    .io_z1(Swapper_508_io_z1)
  );
  Swapper Swapper_509 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_509_io_a0),
    .io_a1(Swapper_509_io_a1),
    .io_z0(Swapper_509_io_z0),
    .io_z1(Swapper_509_io_z1)
  );
  Swapper Swapper_510 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_510_io_a0),
    .io_a1(Swapper_510_io_a1),
    .io_z0(Swapper_510_io_z0),
    .io_z1(Swapper_510_io_z1)
  );
  Swapper Swapper_511 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_511_io_a0),
    .io_a1(Swapper_511_io_a1),
    .io_z0(Swapper_511_io_z0),
    .io_z1(Swapper_511_io_z1)
  );
  Swapper Swapper_512 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_512_io_a0),
    .io_a1(Swapper_512_io_a1),
    .io_z0(Swapper_512_io_z0),
    .io_z1(Swapper_512_io_z1)
  );
  Swapper Swapper_513 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_513_io_a0),
    .io_a1(Swapper_513_io_a1),
    .io_z0(Swapper_513_io_z0),
    .io_z1(Swapper_513_io_z1)
  );
  Swapper Swapper_514 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_514_io_a0),
    .io_a1(Swapper_514_io_a1),
    .io_z0(Swapper_514_io_z0),
    .io_z1(Swapper_514_io_z1)
  );
  Swapper Swapper_515 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_515_io_a0),
    .io_a1(Swapper_515_io_a1),
    .io_z0(Swapper_515_io_z0),
    .io_z1(Swapper_515_io_z1)
  );
  Swapper Swapper_516 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_516_io_a0),
    .io_a1(Swapper_516_io_a1),
    .io_z0(Swapper_516_io_z0),
    .io_z1(Swapper_516_io_z1)
  );
  Swapper Swapper_517 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_517_io_a0),
    .io_a1(Swapper_517_io_a1),
    .io_z0(Swapper_517_io_z0),
    .io_z1(Swapper_517_io_z1)
  );
  Swapper Swapper_518 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_518_io_a0),
    .io_a1(Swapper_518_io_a1),
    .io_z0(Swapper_518_io_z0),
    .io_z1(Swapper_518_io_z1)
  );
  Swapper Swapper_519 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_519_io_a0),
    .io_a1(Swapper_519_io_a1),
    .io_z0(Swapper_519_io_z0),
    .io_z1(Swapper_519_io_z1)
  );
  Swapper Swapper_520 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_520_io_a0),
    .io_a1(Swapper_520_io_a1),
    .io_z0(Swapper_520_io_z0),
    .io_z1(Swapper_520_io_z1)
  );
  Swapper Swapper_521 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_521_io_a0),
    .io_a1(Swapper_521_io_a1),
    .io_z0(Swapper_521_io_z0),
    .io_z1(Swapper_521_io_z1)
  );
  Swapper Swapper_522 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_522_io_a0),
    .io_a1(Swapper_522_io_a1),
    .io_z0(Swapper_522_io_z0),
    .io_z1(Swapper_522_io_z1)
  );
  Swapper Swapper_523 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_523_io_a0),
    .io_a1(Swapper_523_io_a1),
    .io_z0(Swapper_523_io_z0),
    .io_z1(Swapper_523_io_z1)
  );
  Swapper Swapper_524 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_524_io_a0),
    .io_a1(Swapper_524_io_a1),
    .io_z0(Swapper_524_io_z0),
    .io_z1(Swapper_524_io_z1)
  );
  Swapper Swapper_525 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_525_io_a0),
    .io_a1(Swapper_525_io_a1),
    .io_z0(Swapper_525_io_z0),
    .io_z1(Swapper_525_io_z1)
  );
  Swapper Swapper_526 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_526_io_a0),
    .io_a1(Swapper_526_io_a1),
    .io_z0(Swapper_526_io_z0),
    .io_z1(Swapper_526_io_z1)
  );
  Swapper Swapper_527 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_527_io_a0),
    .io_a1(Swapper_527_io_a1),
    .io_z0(Swapper_527_io_z0),
    .io_z1(Swapper_527_io_z1)
  );
  Swapper Swapper_528 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_528_io_a0),
    .io_a1(Swapper_528_io_a1),
    .io_z0(Swapper_528_io_z0),
    .io_z1(Swapper_528_io_z1)
  );
  Swapper Swapper_529 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_529_io_a0),
    .io_a1(Swapper_529_io_a1),
    .io_z0(Swapper_529_io_z0),
    .io_z1(Swapper_529_io_z1)
  );
  Swapper Swapper_530 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_530_io_a0),
    .io_a1(Swapper_530_io_a1),
    .io_z0(Swapper_530_io_z0),
    .io_z1(Swapper_530_io_z1)
  );
  Swapper Swapper_531 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_531_io_a0),
    .io_a1(Swapper_531_io_a1),
    .io_z0(Swapper_531_io_z0),
    .io_z1(Swapper_531_io_z1)
  );
  Swapper Swapper_532 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_532_io_a0),
    .io_a1(Swapper_532_io_a1),
    .io_z0(Swapper_532_io_z0),
    .io_z1(Swapper_532_io_z1)
  );
  Swapper Swapper_533 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_533_io_a0),
    .io_a1(Swapper_533_io_a1),
    .io_z0(Swapper_533_io_z0),
    .io_z1(Swapper_533_io_z1)
  );
  Swapper Swapper_534 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_534_io_a0),
    .io_a1(Swapper_534_io_a1),
    .io_z0(Swapper_534_io_z0),
    .io_z1(Swapper_534_io_z1)
  );
  Swapper Swapper_535 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_535_io_a0),
    .io_a1(Swapper_535_io_a1),
    .io_z0(Swapper_535_io_z0),
    .io_z1(Swapper_535_io_z1)
  );
  Swapper Swapper_536 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_536_io_a0),
    .io_a1(Swapper_536_io_a1),
    .io_z0(Swapper_536_io_z0),
    .io_z1(Swapper_536_io_z1)
  );
  Swapper Swapper_537 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_537_io_a0),
    .io_a1(Swapper_537_io_a1),
    .io_z0(Swapper_537_io_z0),
    .io_z1(Swapper_537_io_z1)
  );
  Swapper Swapper_538 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_538_io_a0),
    .io_a1(Swapper_538_io_a1),
    .io_z0(Swapper_538_io_z0),
    .io_z1(Swapper_538_io_z1)
  );
  Swapper Swapper_539 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_539_io_a0),
    .io_a1(Swapper_539_io_a1),
    .io_z0(Swapper_539_io_z0),
    .io_z1(Swapper_539_io_z1)
  );
  Swapper Swapper_540 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_540_io_a0),
    .io_a1(Swapper_540_io_a1),
    .io_z0(Swapper_540_io_z0),
    .io_z1(Swapper_540_io_z1)
  );
  Swapper Swapper_541 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_541_io_a0),
    .io_a1(Swapper_541_io_a1),
    .io_z0(Swapper_541_io_z0),
    .io_z1(Swapper_541_io_z1)
  );
  Swapper Swapper_542 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_542_io_a0),
    .io_a1(Swapper_542_io_a1),
    .io_z0(Swapper_542_io_z0),
    .io_z1(Swapper_542_io_z1)
  );
  Swapper Swapper_543 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_543_io_a0),
    .io_a1(Swapper_543_io_a1),
    .io_z0(Swapper_543_io_z0),
    .io_z1(Swapper_543_io_z1)
  );
  Swapper Swapper_544 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_544_io_a0),
    .io_a1(Swapper_544_io_a1),
    .io_z0(Swapper_544_io_z0),
    .io_z1(Swapper_544_io_z1)
  );
  Swapper Swapper_545 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_545_io_a0),
    .io_a1(Swapper_545_io_a1),
    .io_z0(Swapper_545_io_z0),
    .io_z1(Swapper_545_io_z1)
  );
  Swapper Swapper_546 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_546_io_a0),
    .io_a1(Swapper_546_io_a1),
    .io_z0(Swapper_546_io_z0),
    .io_z1(Swapper_546_io_z1)
  );
  Swapper Swapper_547 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_547_io_a0),
    .io_a1(Swapper_547_io_a1),
    .io_z0(Swapper_547_io_z0),
    .io_z1(Swapper_547_io_z1)
  );
  Swapper Swapper_548 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_548_io_a0),
    .io_a1(Swapper_548_io_a1),
    .io_z0(Swapper_548_io_z0),
    .io_z1(Swapper_548_io_z1)
  );
  Swapper Swapper_549 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_549_io_a0),
    .io_a1(Swapper_549_io_a1),
    .io_z0(Swapper_549_io_z0),
    .io_z1(Swapper_549_io_z1)
  );
  Swapper Swapper_550 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_550_io_a0),
    .io_a1(Swapper_550_io_a1),
    .io_z0(Swapper_550_io_z0),
    .io_z1(Swapper_550_io_z1)
  );
  Swapper Swapper_551 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_551_io_a0),
    .io_a1(Swapper_551_io_a1),
    .io_z0(Swapper_551_io_z0),
    .io_z1(Swapper_551_io_z1)
  );
  Swapper Swapper_552 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_552_io_a0),
    .io_a1(Swapper_552_io_a1),
    .io_z0(Swapper_552_io_z0),
    .io_z1(Swapper_552_io_z1)
  );
  Swapper Swapper_553 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_553_io_a0),
    .io_a1(Swapper_553_io_a1),
    .io_z0(Swapper_553_io_z0),
    .io_z1(Swapper_553_io_z1)
  );
  Swapper Swapper_554 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_554_io_a0),
    .io_a1(Swapper_554_io_a1),
    .io_z0(Swapper_554_io_z0),
    .io_z1(Swapper_554_io_z1)
  );
  Swapper Swapper_555 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_555_io_a0),
    .io_a1(Swapper_555_io_a1),
    .io_z0(Swapper_555_io_z0),
    .io_z1(Swapper_555_io_z1)
  );
  Swapper Swapper_556 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_556_io_a0),
    .io_a1(Swapper_556_io_a1),
    .io_z0(Swapper_556_io_z0),
    .io_z1(Swapper_556_io_z1)
  );
  Swapper Swapper_557 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_557_io_a0),
    .io_a1(Swapper_557_io_a1),
    .io_z0(Swapper_557_io_z0),
    .io_z1(Swapper_557_io_z1)
  );
  Swapper Swapper_558 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_558_io_a0),
    .io_a1(Swapper_558_io_a1),
    .io_z0(Swapper_558_io_z0),
    .io_z1(Swapper_558_io_z1)
  );
  Swapper Swapper_559 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_559_io_a0),
    .io_a1(Swapper_559_io_a1),
    .io_z0(Swapper_559_io_z0),
    .io_z1(Swapper_559_io_z1)
  );
  Swapper Swapper_560 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_560_io_a0),
    .io_a1(Swapper_560_io_a1),
    .io_z0(Swapper_560_io_z0),
    .io_z1(Swapper_560_io_z1)
  );
  Swapper Swapper_561 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_561_io_a0),
    .io_a1(Swapper_561_io_a1),
    .io_z0(Swapper_561_io_z0),
    .io_z1(Swapper_561_io_z1)
  );
  Swapper Swapper_562 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_562_io_a0),
    .io_a1(Swapper_562_io_a1),
    .io_z0(Swapper_562_io_z0),
    .io_z1(Swapper_562_io_z1)
  );
  Swapper Swapper_563 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_563_io_a0),
    .io_a1(Swapper_563_io_a1),
    .io_z0(Swapper_563_io_z0),
    .io_z1(Swapper_563_io_z1)
  );
  Swapper Swapper_564 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_564_io_a0),
    .io_a1(Swapper_564_io_a1),
    .io_z0(Swapper_564_io_z0),
    .io_z1(Swapper_564_io_z1)
  );
  Swapper Swapper_565 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_565_io_a0),
    .io_a1(Swapper_565_io_a1),
    .io_z0(Swapper_565_io_z0),
    .io_z1(Swapper_565_io_z1)
  );
  Swapper Swapper_566 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_566_io_a0),
    .io_a1(Swapper_566_io_a1),
    .io_z0(Swapper_566_io_z0),
    .io_z1(Swapper_566_io_z1)
  );
  Swapper Swapper_567 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_567_io_a0),
    .io_a1(Swapper_567_io_a1),
    .io_z0(Swapper_567_io_z0),
    .io_z1(Swapper_567_io_z1)
  );
  Swapper Swapper_568 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_568_io_a0),
    .io_a1(Swapper_568_io_a1),
    .io_z0(Swapper_568_io_z0),
    .io_z1(Swapper_568_io_z1)
  );
  Swapper Swapper_569 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_569_io_a0),
    .io_a1(Swapper_569_io_a1),
    .io_z0(Swapper_569_io_z0),
    .io_z1(Swapper_569_io_z1)
  );
  Swapper Swapper_570 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_570_io_a0),
    .io_a1(Swapper_570_io_a1),
    .io_z0(Swapper_570_io_z0),
    .io_z1(Swapper_570_io_z1)
  );
  Swapper Swapper_571 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_571_io_a0),
    .io_a1(Swapper_571_io_a1),
    .io_z0(Swapper_571_io_z0),
    .io_z1(Swapper_571_io_z1)
  );
  Swapper Swapper_572 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_572_io_a0),
    .io_a1(Swapper_572_io_a1),
    .io_z0(Swapper_572_io_z0),
    .io_z1(Swapper_572_io_z1)
  );
  Swapper Swapper_573 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_573_io_a0),
    .io_a1(Swapper_573_io_a1),
    .io_z0(Swapper_573_io_z0),
    .io_z1(Swapper_573_io_z1)
  );
  Swapper Swapper_574 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_574_io_a0),
    .io_a1(Swapper_574_io_a1),
    .io_z0(Swapper_574_io_z0),
    .io_z1(Swapper_574_io_z1)
  );
  Swapper Swapper_575 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_575_io_a0),
    .io_a1(Swapper_575_io_a1),
    .io_z0(Swapper_575_io_z0),
    .io_z1(Swapper_575_io_z1)
  );
  Swapper Swapper_576 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_576_io_a0),
    .io_a1(Swapper_576_io_a1),
    .io_z0(Swapper_576_io_z0),
    .io_z1(Swapper_576_io_z1)
  );
  Swapper Swapper_577 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_577_io_a0),
    .io_a1(Swapper_577_io_a1),
    .io_z0(Swapper_577_io_z0),
    .io_z1(Swapper_577_io_z1)
  );
  Swapper Swapper_578 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_578_io_a0),
    .io_a1(Swapper_578_io_a1),
    .io_z0(Swapper_578_io_z0),
    .io_z1(Swapper_578_io_z1)
  );
  Swapper Swapper_579 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_579_io_a0),
    .io_a1(Swapper_579_io_a1),
    .io_z0(Swapper_579_io_z0),
    .io_z1(Swapper_579_io_z1)
  );
  Swapper Swapper_580 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_580_io_a0),
    .io_a1(Swapper_580_io_a1),
    .io_z0(Swapper_580_io_z0),
    .io_z1(Swapper_580_io_z1)
  );
  Swapper Swapper_581 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_581_io_a0),
    .io_a1(Swapper_581_io_a1),
    .io_z0(Swapper_581_io_z0),
    .io_z1(Swapper_581_io_z1)
  );
  Swapper Swapper_582 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_582_io_a0),
    .io_a1(Swapper_582_io_a1),
    .io_z0(Swapper_582_io_z0),
    .io_z1(Swapper_582_io_z1)
  );
  Swapper Swapper_583 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_583_io_a0),
    .io_a1(Swapper_583_io_a1),
    .io_z0(Swapper_583_io_z0),
    .io_z1(Swapper_583_io_z1)
  );
  Swapper Swapper_584 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_584_io_a0),
    .io_a1(Swapper_584_io_a1),
    .io_z0(Swapper_584_io_z0),
    .io_z1(Swapper_584_io_z1)
  );
  Swapper Swapper_585 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_585_io_a0),
    .io_a1(Swapper_585_io_a1),
    .io_z0(Swapper_585_io_z0),
    .io_z1(Swapper_585_io_z1)
  );
  Swapper Swapper_586 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_586_io_a0),
    .io_a1(Swapper_586_io_a1),
    .io_z0(Swapper_586_io_z0),
    .io_z1(Swapper_586_io_z1)
  );
  Swapper Swapper_587 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_587_io_a0),
    .io_a1(Swapper_587_io_a1),
    .io_z0(Swapper_587_io_z0),
    .io_z1(Swapper_587_io_z1)
  );
  Swapper Swapper_588 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_588_io_a0),
    .io_a1(Swapper_588_io_a1),
    .io_z0(Swapper_588_io_z0),
    .io_z1(Swapper_588_io_z1)
  );
  Swapper Swapper_589 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_589_io_a0),
    .io_a1(Swapper_589_io_a1),
    .io_z0(Swapper_589_io_z0),
    .io_z1(Swapper_589_io_z1)
  );
  Swapper Swapper_590 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_590_io_a0),
    .io_a1(Swapper_590_io_a1),
    .io_z0(Swapper_590_io_z0),
    .io_z1(Swapper_590_io_z1)
  );
  Swapper Swapper_591 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_591_io_a0),
    .io_a1(Swapper_591_io_a1),
    .io_z0(Swapper_591_io_z0),
    .io_z1(Swapper_591_io_z1)
  );
  Swapper Swapper_592 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_592_io_a0),
    .io_a1(Swapper_592_io_a1),
    .io_z0(Swapper_592_io_z0),
    .io_z1(Swapper_592_io_z1)
  );
  Swapper Swapper_593 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_593_io_a0),
    .io_a1(Swapper_593_io_a1),
    .io_z0(Swapper_593_io_z0),
    .io_z1(Swapper_593_io_z1)
  );
  Swapper Swapper_594 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_594_io_a0),
    .io_a1(Swapper_594_io_a1),
    .io_z0(Swapper_594_io_z0),
    .io_z1(Swapper_594_io_z1)
  );
  Swapper Swapper_595 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_595_io_a0),
    .io_a1(Swapper_595_io_a1),
    .io_z0(Swapper_595_io_z0),
    .io_z1(Swapper_595_io_z1)
  );
  Swapper Swapper_596 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_596_io_a0),
    .io_a1(Swapper_596_io_a1),
    .io_z0(Swapper_596_io_z0),
    .io_z1(Swapper_596_io_z1)
  );
  Swapper Swapper_597 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_597_io_a0),
    .io_a1(Swapper_597_io_a1),
    .io_z0(Swapper_597_io_z0),
    .io_z1(Swapper_597_io_z1)
  );
  Swapper Swapper_598 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_598_io_a0),
    .io_a1(Swapper_598_io_a1),
    .io_z0(Swapper_598_io_z0),
    .io_z1(Swapper_598_io_z1)
  );
  Swapper Swapper_599 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_599_io_a0),
    .io_a1(Swapper_599_io_a1),
    .io_z0(Swapper_599_io_z0),
    .io_z1(Swapper_599_io_z1)
  );
  Swapper Swapper_600 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_600_io_a0),
    .io_a1(Swapper_600_io_a1),
    .io_z0(Swapper_600_io_z0),
    .io_z1(Swapper_600_io_z1)
  );
  Swapper Swapper_601 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_601_io_a0),
    .io_a1(Swapper_601_io_a1),
    .io_z0(Swapper_601_io_z0),
    .io_z1(Swapper_601_io_z1)
  );
  Swapper Swapper_602 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_602_io_a0),
    .io_a1(Swapper_602_io_a1),
    .io_z0(Swapper_602_io_z0),
    .io_z1(Swapper_602_io_z1)
  );
  Swapper Swapper_603 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_603_io_a0),
    .io_a1(Swapper_603_io_a1),
    .io_z0(Swapper_603_io_z0),
    .io_z1(Swapper_603_io_z1)
  );
  Swapper Swapper_604 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_604_io_a0),
    .io_a1(Swapper_604_io_a1),
    .io_z0(Swapper_604_io_z0),
    .io_z1(Swapper_604_io_z1)
  );
  Swapper Swapper_605 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_605_io_a0),
    .io_a1(Swapper_605_io_a1),
    .io_z0(Swapper_605_io_z0),
    .io_z1(Swapper_605_io_z1)
  );
  Swapper Swapper_606 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_606_io_a0),
    .io_a1(Swapper_606_io_a1),
    .io_z0(Swapper_606_io_z0),
    .io_z1(Swapper_606_io_z1)
  );
  Swapper Swapper_607 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_607_io_a0),
    .io_a1(Swapper_607_io_a1),
    .io_z0(Swapper_607_io_z0),
    .io_z1(Swapper_607_io_z1)
  );
  Swapper Swapper_608 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_608_io_a0),
    .io_a1(Swapper_608_io_a1),
    .io_z0(Swapper_608_io_z0),
    .io_z1(Swapper_608_io_z1)
  );
  Swapper Swapper_609 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_609_io_a0),
    .io_a1(Swapper_609_io_a1),
    .io_z0(Swapper_609_io_z0),
    .io_z1(Swapper_609_io_z1)
  );
  Swapper Swapper_610 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_610_io_a0),
    .io_a1(Swapper_610_io_a1),
    .io_z0(Swapper_610_io_z0),
    .io_z1(Swapper_610_io_z1)
  );
  Swapper Swapper_611 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_611_io_a0),
    .io_a1(Swapper_611_io_a1),
    .io_z0(Swapper_611_io_z0),
    .io_z1(Swapper_611_io_z1)
  );
  Swapper Swapper_612 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_612_io_a0),
    .io_a1(Swapper_612_io_a1),
    .io_z0(Swapper_612_io_z0),
    .io_z1(Swapper_612_io_z1)
  );
  Swapper Swapper_613 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_613_io_a0),
    .io_a1(Swapper_613_io_a1),
    .io_z0(Swapper_613_io_z0),
    .io_z1(Swapper_613_io_z1)
  );
  Swapper Swapper_614 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_614_io_a0),
    .io_a1(Swapper_614_io_a1),
    .io_z0(Swapper_614_io_z0),
    .io_z1(Swapper_614_io_z1)
  );
  Swapper Swapper_615 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_615_io_a0),
    .io_a1(Swapper_615_io_a1),
    .io_z0(Swapper_615_io_z0),
    .io_z1(Swapper_615_io_z1)
  );
  Swapper Swapper_616 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_616_io_a0),
    .io_a1(Swapper_616_io_a1),
    .io_z0(Swapper_616_io_z0),
    .io_z1(Swapper_616_io_z1)
  );
  Swapper Swapper_617 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_617_io_a0),
    .io_a1(Swapper_617_io_a1),
    .io_z0(Swapper_617_io_z0),
    .io_z1(Swapper_617_io_z1)
  );
  Swapper Swapper_618 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_618_io_a0),
    .io_a1(Swapper_618_io_a1),
    .io_z0(Swapper_618_io_z0),
    .io_z1(Swapper_618_io_z1)
  );
  Swapper Swapper_619 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_619_io_a0),
    .io_a1(Swapper_619_io_a1),
    .io_z0(Swapper_619_io_z0),
    .io_z1(Swapper_619_io_z1)
  );
  Swapper Swapper_620 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_620_io_a0),
    .io_a1(Swapper_620_io_a1),
    .io_z0(Swapper_620_io_z0),
    .io_z1(Swapper_620_io_z1)
  );
  Swapper Swapper_621 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_621_io_a0),
    .io_a1(Swapper_621_io_a1),
    .io_z0(Swapper_621_io_z0),
    .io_z1(Swapper_621_io_z1)
  );
  Swapper Swapper_622 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_622_io_a0),
    .io_a1(Swapper_622_io_a1),
    .io_z0(Swapper_622_io_z0),
    .io_z1(Swapper_622_io_z1)
  );
  Swapper Swapper_623 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_623_io_a0),
    .io_a1(Swapper_623_io_a1),
    .io_z0(Swapper_623_io_z0),
    .io_z1(Swapper_623_io_z1)
  );
  Swapper Swapper_624 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_624_io_a0),
    .io_a1(Swapper_624_io_a1),
    .io_z0(Swapper_624_io_z0),
    .io_z1(Swapper_624_io_z1)
  );
  Swapper Swapper_625 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_625_io_a0),
    .io_a1(Swapper_625_io_a1),
    .io_z0(Swapper_625_io_z0),
    .io_z1(Swapper_625_io_z1)
  );
  Swapper Swapper_626 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_626_io_a0),
    .io_a1(Swapper_626_io_a1),
    .io_z0(Swapper_626_io_z0),
    .io_z1(Swapper_626_io_z1)
  );
  Swapper Swapper_627 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_627_io_a0),
    .io_a1(Swapper_627_io_a1),
    .io_z0(Swapper_627_io_z0),
    .io_z1(Swapper_627_io_z1)
  );
  Swapper Swapper_628 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_628_io_a0),
    .io_a1(Swapper_628_io_a1),
    .io_z0(Swapper_628_io_z0),
    .io_z1(Swapper_628_io_z1)
  );
  Swapper Swapper_629 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_629_io_a0),
    .io_a1(Swapper_629_io_a1),
    .io_z0(Swapper_629_io_z0),
    .io_z1(Swapper_629_io_z1)
  );
  Swapper Swapper_630 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_630_io_a0),
    .io_a1(Swapper_630_io_a1),
    .io_z0(Swapper_630_io_z0),
    .io_z1(Swapper_630_io_z1)
  );
  Swapper Swapper_631 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_631_io_a0),
    .io_a1(Swapper_631_io_a1),
    .io_z0(Swapper_631_io_z0),
    .io_z1(Swapper_631_io_z1)
  );
  Swapper Swapper_632 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_632_io_a0),
    .io_a1(Swapper_632_io_a1),
    .io_z0(Swapper_632_io_z0),
    .io_z1(Swapper_632_io_z1)
  );
  Swapper Swapper_633 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_633_io_a0),
    .io_a1(Swapper_633_io_a1),
    .io_z0(Swapper_633_io_z0),
    .io_z1(Swapper_633_io_z1)
  );
  Swapper Swapper_634 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_634_io_a0),
    .io_a1(Swapper_634_io_a1),
    .io_z0(Swapper_634_io_z0),
    .io_z1(Swapper_634_io_z1)
  );
  Swapper Swapper_635 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_635_io_a0),
    .io_a1(Swapper_635_io_a1),
    .io_z0(Swapper_635_io_z0),
    .io_z1(Swapper_635_io_z1)
  );
  Swapper Swapper_636 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_636_io_a0),
    .io_a1(Swapper_636_io_a1),
    .io_z0(Swapper_636_io_z0),
    .io_z1(Swapper_636_io_z1)
  );
  Swapper Swapper_637 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_637_io_a0),
    .io_a1(Swapper_637_io_a1),
    .io_z0(Swapper_637_io_z0),
    .io_z1(Swapper_637_io_z1)
  );
  Swapper Swapper_638 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_638_io_a0),
    .io_a1(Swapper_638_io_a1),
    .io_z0(Swapper_638_io_z0),
    .io_z1(Swapper_638_io_z1)
  );
  Swapper Swapper_639 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_639_io_a0),
    .io_a1(Swapper_639_io_a1),
    .io_z0(Swapper_639_io_z0),
    .io_z1(Swapper_639_io_z1)
  );
  Swapper Swapper_640 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_640_io_a0),
    .io_a1(Swapper_640_io_a1),
    .io_z0(Swapper_640_io_z0),
    .io_z1(Swapper_640_io_z1)
  );
  Swapper Swapper_641 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_641_io_a0),
    .io_a1(Swapper_641_io_a1),
    .io_z0(Swapper_641_io_z0),
    .io_z1(Swapper_641_io_z1)
  );
  Swapper Swapper_642 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_642_io_a0),
    .io_a1(Swapper_642_io_a1),
    .io_z0(Swapper_642_io_z0),
    .io_z1(Swapper_642_io_z1)
  );
  Swapper Swapper_643 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_643_io_a0),
    .io_a1(Swapper_643_io_a1),
    .io_z0(Swapper_643_io_z0),
    .io_z1(Swapper_643_io_z1)
  );
  Swapper Swapper_644 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_644_io_a0),
    .io_a1(Swapper_644_io_a1),
    .io_z0(Swapper_644_io_z0),
    .io_z1(Swapper_644_io_z1)
  );
  Swapper Swapper_645 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_645_io_a0),
    .io_a1(Swapper_645_io_a1),
    .io_z0(Swapper_645_io_z0),
    .io_z1(Swapper_645_io_z1)
  );
  Swapper Swapper_646 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_646_io_a0),
    .io_a1(Swapper_646_io_a1),
    .io_z0(Swapper_646_io_z0),
    .io_z1(Swapper_646_io_z1)
  );
  Swapper Swapper_647 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_647_io_a0),
    .io_a1(Swapper_647_io_a1),
    .io_z0(Swapper_647_io_z0),
    .io_z1(Swapper_647_io_z1)
  );
  Swapper Swapper_648 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_648_io_a0),
    .io_a1(Swapper_648_io_a1),
    .io_z0(Swapper_648_io_z0),
    .io_z1(Swapper_648_io_z1)
  );
  Swapper Swapper_649 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_649_io_a0),
    .io_a1(Swapper_649_io_a1),
    .io_z0(Swapper_649_io_z0),
    .io_z1(Swapper_649_io_z1)
  );
  Swapper Swapper_650 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_650_io_a0),
    .io_a1(Swapper_650_io_a1),
    .io_z0(Swapper_650_io_z0),
    .io_z1(Swapper_650_io_z1)
  );
  Swapper Swapper_651 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_651_io_a0),
    .io_a1(Swapper_651_io_a1),
    .io_z0(Swapper_651_io_z0),
    .io_z1(Swapper_651_io_z1)
  );
  Swapper Swapper_652 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_652_io_a0),
    .io_a1(Swapper_652_io_a1),
    .io_z0(Swapper_652_io_z0),
    .io_z1(Swapper_652_io_z1)
  );
  Swapper Swapper_653 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_653_io_a0),
    .io_a1(Swapper_653_io_a1),
    .io_z0(Swapper_653_io_z0),
    .io_z1(Swapper_653_io_z1)
  );
  Swapper Swapper_654 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_654_io_a0),
    .io_a1(Swapper_654_io_a1),
    .io_z0(Swapper_654_io_z0),
    .io_z1(Swapper_654_io_z1)
  );
  Swapper Swapper_655 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_655_io_a0),
    .io_a1(Swapper_655_io_a1),
    .io_z0(Swapper_655_io_z0),
    .io_z1(Swapper_655_io_z1)
  );
  Swapper Swapper_656 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_656_io_a0),
    .io_a1(Swapper_656_io_a1),
    .io_z0(Swapper_656_io_z0),
    .io_z1(Swapper_656_io_z1)
  );
  Swapper Swapper_657 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_657_io_a0),
    .io_a1(Swapper_657_io_a1),
    .io_z0(Swapper_657_io_z0),
    .io_z1(Swapper_657_io_z1)
  );
  Swapper Swapper_658 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_658_io_a0),
    .io_a1(Swapper_658_io_a1),
    .io_z0(Swapper_658_io_z0),
    .io_z1(Swapper_658_io_z1)
  );
  Swapper Swapper_659 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_659_io_a0),
    .io_a1(Swapper_659_io_a1),
    .io_z0(Swapper_659_io_z0),
    .io_z1(Swapper_659_io_z1)
  );
  Swapper Swapper_660 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_660_io_a0),
    .io_a1(Swapper_660_io_a1),
    .io_z0(Swapper_660_io_z0),
    .io_z1(Swapper_660_io_z1)
  );
  Swapper Swapper_661 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_661_io_a0),
    .io_a1(Swapper_661_io_a1),
    .io_z0(Swapper_661_io_z0),
    .io_z1(Swapper_661_io_z1)
  );
  Swapper Swapper_662 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_662_io_a0),
    .io_a1(Swapper_662_io_a1),
    .io_z0(Swapper_662_io_z0),
    .io_z1(Swapper_662_io_z1)
  );
  Swapper Swapper_663 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_663_io_a0),
    .io_a1(Swapper_663_io_a1),
    .io_z0(Swapper_663_io_z0),
    .io_z1(Swapper_663_io_z1)
  );
  Swapper Swapper_664 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_664_io_a0),
    .io_a1(Swapper_664_io_a1),
    .io_z0(Swapper_664_io_z0),
    .io_z1(Swapper_664_io_z1)
  );
  Swapper Swapper_665 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_665_io_a0),
    .io_a1(Swapper_665_io_a1),
    .io_z0(Swapper_665_io_z0),
    .io_z1(Swapper_665_io_z1)
  );
  Swapper Swapper_666 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_666_io_a0),
    .io_a1(Swapper_666_io_a1),
    .io_z0(Swapper_666_io_z0),
    .io_z1(Swapper_666_io_z1)
  );
  Swapper Swapper_667 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_667_io_a0),
    .io_a1(Swapper_667_io_a1),
    .io_z0(Swapper_667_io_z0),
    .io_z1(Swapper_667_io_z1)
  );
  Swapper Swapper_668 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_668_io_a0),
    .io_a1(Swapper_668_io_a1),
    .io_z0(Swapper_668_io_z0),
    .io_z1(Swapper_668_io_z1)
  );
  Swapper Swapper_669 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_669_io_a0),
    .io_a1(Swapper_669_io_a1),
    .io_z0(Swapper_669_io_z0),
    .io_z1(Swapper_669_io_z1)
  );
  Swapper Swapper_670 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_670_io_a0),
    .io_a1(Swapper_670_io_a1),
    .io_z0(Swapper_670_io_z0),
    .io_z1(Swapper_670_io_z1)
  );
  Swapper Swapper_671 ( // @[bitonic_sort.scala 31:25]
    .io_a0(Swapper_671_io_a0),
    .io_a1(Swapper_671_io_a1),
    .io_z0(Swapper_671_io_z0),
    .io_z1(Swapper_671_io_z1)
  );
  assign io_z_0 = Swapper_640_io_z0; // @[bitonic_sort.scala 58:8]
  assign io_z_1 = Swapper_640_io_z1; // @[bitonic_sort.scala 58:8]
  assign io_z_2 = Swapper_641_io_z0; // @[bitonic_sort.scala 58:8]
  assign io_z_3 = Swapper_641_io_z1; // @[bitonic_sort.scala 58:8]
  assign io_z_4 = Swapper_642_io_z0; // @[bitonic_sort.scala 58:8]
  assign io_z_5 = Swapper_642_io_z1; // @[bitonic_sort.scala 58:8]
  assign io_z_6 = Swapper_643_io_z0; // @[bitonic_sort.scala 58:8]
  assign io_z_7 = Swapper_643_io_z1; // @[bitonic_sort.scala 58:8]
  assign io_z_8 = Swapper_644_io_z0; // @[bitonic_sort.scala 58:8]
  assign io_z_9 = Swapper_644_io_z1; // @[bitonic_sort.scala 58:8]
  assign io_z_10 = Swapper_645_io_z0; // @[bitonic_sort.scala 58:8]
  assign io_z_11 = Swapper_645_io_z1; // @[bitonic_sort.scala 58:8]
  assign io_z_12 = Swapper_646_io_z0; // @[bitonic_sort.scala 58:8]
  assign io_z_13 = Swapper_646_io_z1; // @[bitonic_sort.scala 58:8]
  assign io_z_14 = Swapper_647_io_z0; // @[bitonic_sort.scala 58:8]
  assign io_z_15 = Swapper_647_io_z1; // @[bitonic_sort.scala 58:8]
  assign io_z_16 = Swapper_648_io_z0; // @[bitonic_sort.scala 58:8]
  assign io_z_17 = Swapper_648_io_z1; // @[bitonic_sort.scala 58:8]
  assign io_z_18 = Swapper_649_io_z0; // @[bitonic_sort.scala 58:8]
  assign io_z_19 = Swapper_649_io_z1; // @[bitonic_sort.scala 58:8]
  assign io_z_20 = Swapper_650_io_z0; // @[bitonic_sort.scala 58:8]
  assign io_z_21 = Swapper_650_io_z1; // @[bitonic_sort.scala 58:8]
  assign io_z_22 = Swapper_651_io_z0; // @[bitonic_sort.scala 58:8]
  assign io_z_23 = Swapper_651_io_z1; // @[bitonic_sort.scala 58:8]
  assign io_z_24 = Swapper_652_io_z0; // @[bitonic_sort.scala 58:8]
  assign io_z_25 = Swapper_652_io_z1; // @[bitonic_sort.scala 58:8]
  assign io_z_26 = Swapper_653_io_z0; // @[bitonic_sort.scala 58:8]
  assign io_z_27 = Swapper_653_io_z1; // @[bitonic_sort.scala 58:8]
  assign io_z_28 = Swapper_654_io_z0; // @[bitonic_sort.scala 58:8]
  assign io_z_29 = Swapper_654_io_z1; // @[bitonic_sort.scala 58:8]
  assign io_z_30 = Swapper_655_io_z0; // @[bitonic_sort.scala 58:8]
  assign io_z_31 = Swapper_655_io_z1; // @[bitonic_sort.scala 58:8]
  assign io_z_32 = Swapper_656_io_z0; // @[bitonic_sort.scala 58:8]
  assign io_z_33 = Swapper_656_io_z1; // @[bitonic_sort.scala 58:8]
  assign io_z_34 = Swapper_657_io_z0; // @[bitonic_sort.scala 58:8]
  assign io_z_35 = Swapper_657_io_z1; // @[bitonic_sort.scala 58:8]
  assign io_z_36 = Swapper_658_io_z0; // @[bitonic_sort.scala 58:8]
  assign io_z_37 = Swapper_658_io_z1; // @[bitonic_sort.scala 58:8]
  assign io_z_38 = Swapper_659_io_z0; // @[bitonic_sort.scala 58:8]
  assign io_z_39 = Swapper_659_io_z1; // @[bitonic_sort.scala 58:8]
  assign io_z_40 = Swapper_660_io_z0; // @[bitonic_sort.scala 58:8]
  assign io_z_41 = Swapper_660_io_z1; // @[bitonic_sort.scala 58:8]
  assign io_z_42 = Swapper_661_io_z0; // @[bitonic_sort.scala 58:8]
  assign io_z_43 = Swapper_661_io_z1; // @[bitonic_sort.scala 58:8]
  assign io_z_44 = Swapper_662_io_z0; // @[bitonic_sort.scala 58:8]
  assign io_z_45 = Swapper_662_io_z1; // @[bitonic_sort.scala 58:8]
  assign io_z_46 = Swapper_663_io_z0; // @[bitonic_sort.scala 58:8]
  assign io_z_47 = Swapper_663_io_z1; // @[bitonic_sort.scala 58:8]
  assign io_z_48 = Swapper_664_io_z0; // @[bitonic_sort.scala 58:8]
  assign io_z_49 = Swapper_664_io_z1; // @[bitonic_sort.scala 58:8]
  assign io_z_50 = Swapper_665_io_z0; // @[bitonic_sort.scala 58:8]
  assign io_z_51 = Swapper_665_io_z1; // @[bitonic_sort.scala 58:8]
  assign io_z_52 = Swapper_666_io_z0; // @[bitonic_sort.scala 58:8]
  assign io_z_53 = Swapper_666_io_z1; // @[bitonic_sort.scala 58:8]
  assign io_z_54 = Swapper_667_io_z0; // @[bitonic_sort.scala 58:8]
  assign io_z_55 = Swapper_667_io_z1; // @[bitonic_sort.scala 58:8]
  assign io_z_56 = Swapper_668_io_z0; // @[bitonic_sort.scala 58:8]
  assign io_z_57 = Swapper_668_io_z1; // @[bitonic_sort.scala 58:8]
  assign io_z_58 = Swapper_669_io_z0; // @[bitonic_sort.scala 58:8]
  assign io_z_59 = Swapper_669_io_z1; // @[bitonic_sort.scala 58:8]
  assign io_z_60 = Swapper_670_io_z0; // @[bitonic_sort.scala 58:8]
  assign io_z_61 = Swapper_670_io_z1; // @[bitonic_sort.scala 58:8]
  assign io_z_62 = Swapper_671_io_z0; // @[bitonic_sort.scala 58:8]
  assign io_z_63 = Swapper_671_io_z1; // @[bitonic_sort.scala 58:8]
  assign Swapper_io_a0 = io_a_0; // @[bitonic_sort.scala 32:19]
  assign Swapper_io_a1 = io_a_1; // @[bitonic_sort.scala 33:19]
  assign Swapper_1_io_a0 = io_a_3; // @[bitonic_sort.scala 32:19]
  assign Swapper_1_io_a1 = io_a_2; // @[bitonic_sort.scala 33:19]
  assign Swapper_2_io_a0 = io_a_4; // @[bitonic_sort.scala 32:19]
  assign Swapper_2_io_a1 = io_a_5; // @[bitonic_sort.scala 33:19]
  assign Swapper_3_io_a0 = io_a_7; // @[bitonic_sort.scala 32:19]
  assign Swapper_3_io_a1 = io_a_6; // @[bitonic_sort.scala 33:19]
  assign Swapper_4_io_a0 = io_a_8; // @[bitonic_sort.scala 32:19]
  assign Swapper_4_io_a1 = io_a_9; // @[bitonic_sort.scala 33:19]
  assign Swapper_5_io_a0 = io_a_11; // @[bitonic_sort.scala 32:19]
  assign Swapper_5_io_a1 = io_a_10; // @[bitonic_sort.scala 33:19]
  assign Swapper_6_io_a0 = io_a_12; // @[bitonic_sort.scala 32:19]
  assign Swapper_6_io_a1 = io_a_13; // @[bitonic_sort.scala 33:19]
  assign Swapper_7_io_a0 = io_a_15; // @[bitonic_sort.scala 32:19]
  assign Swapper_7_io_a1 = io_a_14; // @[bitonic_sort.scala 33:19]
  assign Swapper_8_io_a0 = io_a_16; // @[bitonic_sort.scala 32:19]
  assign Swapper_8_io_a1 = io_a_17; // @[bitonic_sort.scala 33:19]
  assign Swapper_9_io_a0 = io_a_19; // @[bitonic_sort.scala 32:19]
  assign Swapper_9_io_a1 = io_a_18; // @[bitonic_sort.scala 33:19]
  assign Swapper_10_io_a0 = io_a_20; // @[bitonic_sort.scala 32:19]
  assign Swapper_10_io_a1 = io_a_21; // @[bitonic_sort.scala 33:19]
  assign Swapper_11_io_a0 = io_a_23; // @[bitonic_sort.scala 32:19]
  assign Swapper_11_io_a1 = io_a_22; // @[bitonic_sort.scala 33:19]
  assign Swapper_12_io_a0 = io_a_24; // @[bitonic_sort.scala 32:19]
  assign Swapper_12_io_a1 = io_a_25; // @[bitonic_sort.scala 33:19]
  assign Swapper_13_io_a0 = io_a_27; // @[bitonic_sort.scala 32:19]
  assign Swapper_13_io_a1 = io_a_26; // @[bitonic_sort.scala 33:19]
  assign Swapper_14_io_a0 = io_a_28; // @[bitonic_sort.scala 32:19]
  assign Swapper_14_io_a1 = io_a_29; // @[bitonic_sort.scala 33:19]
  assign Swapper_15_io_a0 = io_a_31; // @[bitonic_sort.scala 32:19]
  assign Swapper_15_io_a1 = io_a_30; // @[bitonic_sort.scala 33:19]
  assign Swapper_16_io_a0 = io_a_32; // @[bitonic_sort.scala 32:19]
  assign Swapper_16_io_a1 = io_a_33; // @[bitonic_sort.scala 33:19]
  assign Swapper_17_io_a0 = io_a_35; // @[bitonic_sort.scala 32:19]
  assign Swapper_17_io_a1 = io_a_34; // @[bitonic_sort.scala 33:19]
  assign Swapper_18_io_a0 = io_a_36; // @[bitonic_sort.scala 32:19]
  assign Swapper_18_io_a1 = io_a_37; // @[bitonic_sort.scala 33:19]
  assign Swapper_19_io_a0 = io_a_39; // @[bitonic_sort.scala 32:19]
  assign Swapper_19_io_a1 = io_a_38; // @[bitonic_sort.scala 33:19]
  assign Swapper_20_io_a0 = io_a_40; // @[bitonic_sort.scala 32:19]
  assign Swapper_20_io_a1 = io_a_41; // @[bitonic_sort.scala 33:19]
  assign Swapper_21_io_a0 = io_a_43; // @[bitonic_sort.scala 32:19]
  assign Swapper_21_io_a1 = io_a_42; // @[bitonic_sort.scala 33:19]
  assign Swapper_22_io_a0 = io_a_44; // @[bitonic_sort.scala 32:19]
  assign Swapper_22_io_a1 = io_a_45; // @[bitonic_sort.scala 33:19]
  assign Swapper_23_io_a0 = io_a_47; // @[bitonic_sort.scala 32:19]
  assign Swapper_23_io_a1 = io_a_46; // @[bitonic_sort.scala 33:19]
  assign Swapper_24_io_a0 = io_a_48; // @[bitonic_sort.scala 32:19]
  assign Swapper_24_io_a1 = io_a_49; // @[bitonic_sort.scala 33:19]
  assign Swapper_25_io_a0 = io_a_51; // @[bitonic_sort.scala 32:19]
  assign Swapper_25_io_a1 = io_a_50; // @[bitonic_sort.scala 33:19]
  assign Swapper_26_io_a0 = io_a_52; // @[bitonic_sort.scala 32:19]
  assign Swapper_26_io_a1 = io_a_53; // @[bitonic_sort.scala 33:19]
  assign Swapper_27_io_a0 = io_a_55; // @[bitonic_sort.scala 32:19]
  assign Swapper_27_io_a1 = io_a_54; // @[bitonic_sort.scala 33:19]
  assign Swapper_28_io_a0 = io_a_56; // @[bitonic_sort.scala 32:19]
  assign Swapper_28_io_a1 = io_a_57; // @[bitonic_sort.scala 33:19]
  assign Swapper_29_io_a0 = io_a_59; // @[bitonic_sort.scala 32:19]
  assign Swapper_29_io_a1 = io_a_58; // @[bitonic_sort.scala 33:19]
  assign Swapper_30_io_a0 = io_a_60; // @[bitonic_sort.scala 32:19]
  assign Swapper_30_io_a1 = io_a_61; // @[bitonic_sort.scala 33:19]
  assign Swapper_31_io_a0 = io_a_63; // @[bitonic_sort.scala 32:19]
  assign Swapper_31_io_a1 = io_a_62; // @[bitonic_sort.scala 33:19]
  assign Swapper_32_io_a0 = Swapper_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_32_io_a1 = Swapper_1_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_33_io_a0 = Swapper_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_33_io_a1 = Swapper_1_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_34_io_a0 = Swapper_3_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_34_io_a1 = Swapper_2_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_35_io_a0 = Swapper_3_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_35_io_a1 = Swapper_2_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_36_io_a0 = Swapper_4_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_36_io_a1 = Swapper_5_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_37_io_a0 = Swapper_4_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_37_io_a1 = Swapper_5_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_38_io_a0 = Swapper_7_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_38_io_a1 = Swapper_6_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_39_io_a0 = Swapper_7_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_39_io_a1 = Swapper_6_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_40_io_a0 = Swapper_8_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_40_io_a1 = Swapper_9_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_41_io_a0 = Swapper_8_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_41_io_a1 = Swapper_9_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_42_io_a0 = Swapper_11_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_42_io_a1 = Swapper_10_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_43_io_a0 = Swapper_11_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_43_io_a1 = Swapper_10_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_44_io_a0 = Swapper_12_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_44_io_a1 = Swapper_13_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_45_io_a0 = Swapper_12_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_45_io_a1 = Swapper_13_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_46_io_a0 = Swapper_15_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_46_io_a1 = Swapper_14_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_47_io_a0 = Swapper_15_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_47_io_a1 = Swapper_14_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_48_io_a0 = Swapper_16_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_48_io_a1 = Swapper_17_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_49_io_a0 = Swapper_16_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_49_io_a1 = Swapper_17_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_50_io_a0 = Swapper_19_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_50_io_a1 = Swapper_18_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_51_io_a0 = Swapper_19_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_51_io_a1 = Swapper_18_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_52_io_a0 = Swapper_20_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_52_io_a1 = Swapper_21_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_53_io_a0 = Swapper_20_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_53_io_a1 = Swapper_21_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_54_io_a0 = Swapper_23_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_54_io_a1 = Swapper_22_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_55_io_a0 = Swapper_23_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_55_io_a1 = Swapper_22_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_56_io_a0 = Swapper_24_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_56_io_a1 = Swapper_25_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_57_io_a0 = Swapper_24_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_57_io_a1 = Swapper_25_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_58_io_a0 = Swapper_27_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_58_io_a1 = Swapper_26_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_59_io_a0 = Swapper_27_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_59_io_a1 = Swapper_26_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_60_io_a0 = Swapper_28_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_60_io_a1 = Swapper_29_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_61_io_a0 = Swapper_28_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_61_io_a1 = Swapper_29_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_62_io_a0 = Swapper_31_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_62_io_a1 = Swapper_30_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_63_io_a0 = Swapper_31_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_63_io_a1 = Swapper_30_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_64_io_a0 = Swapper_32_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_64_io_a1 = Swapper_33_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_65_io_a0 = Swapper_32_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_65_io_a1 = Swapper_33_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_66_io_a0 = Swapper_35_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_66_io_a1 = Swapper_34_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_67_io_a0 = Swapper_35_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_67_io_a1 = Swapper_34_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_68_io_a0 = Swapper_36_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_68_io_a1 = Swapper_37_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_69_io_a0 = Swapper_36_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_69_io_a1 = Swapper_37_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_70_io_a0 = Swapper_39_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_70_io_a1 = Swapper_38_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_71_io_a0 = Swapper_39_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_71_io_a1 = Swapper_38_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_72_io_a0 = Swapper_40_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_72_io_a1 = Swapper_41_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_73_io_a0 = Swapper_40_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_73_io_a1 = Swapper_41_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_74_io_a0 = Swapper_43_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_74_io_a1 = Swapper_42_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_75_io_a0 = Swapper_43_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_75_io_a1 = Swapper_42_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_76_io_a0 = Swapper_44_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_76_io_a1 = Swapper_45_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_77_io_a0 = Swapper_44_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_77_io_a1 = Swapper_45_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_78_io_a0 = Swapper_47_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_78_io_a1 = Swapper_46_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_79_io_a0 = Swapper_47_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_79_io_a1 = Swapper_46_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_80_io_a0 = Swapper_48_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_80_io_a1 = Swapper_49_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_81_io_a0 = Swapper_48_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_81_io_a1 = Swapper_49_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_82_io_a0 = Swapper_51_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_82_io_a1 = Swapper_50_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_83_io_a0 = Swapper_51_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_83_io_a1 = Swapper_50_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_84_io_a0 = Swapper_52_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_84_io_a1 = Swapper_53_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_85_io_a0 = Swapper_52_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_85_io_a1 = Swapper_53_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_86_io_a0 = Swapper_55_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_86_io_a1 = Swapper_54_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_87_io_a0 = Swapper_55_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_87_io_a1 = Swapper_54_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_88_io_a0 = Swapper_56_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_88_io_a1 = Swapper_57_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_89_io_a0 = Swapper_56_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_89_io_a1 = Swapper_57_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_90_io_a0 = Swapper_59_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_90_io_a1 = Swapper_58_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_91_io_a0 = Swapper_59_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_91_io_a1 = Swapper_58_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_92_io_a0 = Swapper_60_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_92_io_a1 = Swapper_61_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_93_io_a0 = Swapper_60_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_93_io_a1 = Swapper_61_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_94_io_a0 = Swapper_63_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_94_io_a1 = Swapper_62_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_95_io_a0 = Swapper_63_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_95_io_a1 = Swapper_62_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_96_io_a0 = Swapper_64_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_96_io_a1 = Swapper_66_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_97_io_a0 = Swapper_64_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_97_io_a1 = Swapper_66_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_98_io_a0 = Swapper_65_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_98_io_a1 = Swapper_67_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_99_io_a0 = Swapper_65_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_99_io_a1 = Swapper_67_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_100_io_a0 = Swapper_70_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_100_io_a1 = Swapper_68_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_101_io_a0 = Swapper_70_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_101_io_a1 = Swapper_68_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_102_io_a0 = Swapper_71_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_102_io_a1 = Swapper_69_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_103_io_a0 = Swapper_71_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_103_io_a1 = Swapper_69_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_104_io_a0 = Swapper_72_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_104_io_a1 = Swapper_74_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_105_io_a0 = Swapper_72_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_105_io_a1 = Swapper_74_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_106_io_a0 = Swapper_73_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_106_io_a1 = Swapper_75_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_107_io_a0 = Swapper_73_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_107_io_a1 = Swapper_75_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_108_io_a0 = Swapper_78_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_108_io_a1 = Swapper_76_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_109_io_a0 = Swapper_78_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_109_io_a1 = Swapper_76_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_110_io_a0 = Swapper_79_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_110_io_a1 = Swapper_77_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_111_io_a0 = Swapper_79_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_111_io_a1 = Swapper_77_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_112_io_a0 = Swapper_80_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_112_io_a1 = Swapper_82_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_113_io_a0 = Swapper_80_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_113_io_a1 = Swapper_82_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_114_io_a0 = Swapper_81_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_114_io_a1 = Swapper_83_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_115_io_a0 = Swapper_81_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_115_io_a1 = Swapper_83_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_116_io_a0 = Swapper_86_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_116_io_a1 = Swapper_84_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_117_io_a0 = Swapper_86_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_117_io_a1 = Swapper_84_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_118_io_a0 = Swapper_87_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_118_io_a1 = Swapper_85_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_119_io_a0 = Swapper_87_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_119_io_a1 = Swapper_85_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_120_io_a0 = Swapper_88_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_120_io_a1 = Swapper_90_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_121_io_a0 = Swapper_88_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_121_io_a1 = Swapper_90_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_122_io_a0 = Swapper_89_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_122_io_a1 = Swapper_91_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_123_io_a0 = Swapper_89_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_123_io_a1 = Swapper_91_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_124_io_a0 = Swapper_94_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_124_io_a1 = Swapper_92_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_125_io_a0 = Swapper_94_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_125_io_a1 = Swapper_92_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_126_io_a0 = Swapper_95_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_126_io_a1 = Swapper_93_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_127_io_a0 = Swapper_95_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_127_io_a1 = Swapper_93_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_128_io_a0 = Swapper_96_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_128_io_a1 = Swapper_98_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_129_io_a0 = Swapper_97_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_129_io_a1 = Swapper_99_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_130_io_a0 = Swapper_96_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_130_io_a1 = Swapper_98_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_131_io_a0 = Swapper_97_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_131_io_a1 = Swapper_99_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_132_io_a0 = Swapper_102_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_132_io_a1 = Swapper_100_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_133_io_a0 = Swapper_103_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_133_io_a1 = Swapper_101_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_134_io_a0 = Swapper_102_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_134_io_a1 = Swapper_100_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_135_io_a0 = Swapper_103_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_135_io_a1 = Swapper_101_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_136_io_a0 = Swapper_104_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_136_io_a1 = Swapper_106_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_137_io_a0 = Swapper_105_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_137_io_a1 = Swapper_107_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_138_io_a0 = Swapper_104_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_138_io_a1 = Swapper_106_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_139_io_a0 = Swapper_105_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_139_io_a1 = Swapper_107_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_140_io_a0 = Swapper_110_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_140_io_a1 = Swapper_108_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_141_io_a0 = Swapper_111_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_141_io_a1 = Swapper_109_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_142_io_a0 = Swapper_110_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_142_io_a1 = Swapper_108_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_143_io_a0 = Swapper_111_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_143_io_a1 = Swapper_109_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_144_io_a0 = Swapper_112_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_144_io_a1 = Swapper_114_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_145_io_a0 = Swapper_113_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_145_io_a1 = Swapper_115_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_146_io_a0 = Swapper_112_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_146_io_a1 = Swapper_114_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_147_io_a0 = Swapper_113_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_147_io_a1 = Swapper_115_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_148_io_a0 = Swapper_118_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_148_io_a1 = Swapper_116_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_149_io_a0 = Swapper_119_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_149_io_a1 = Swapper_117_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_150_io_a0 = Swapper_118_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_150_io_a1 = Swapper_116_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_151_io_a0 = Swapper_119_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_151_io_a1 = Swapper_117_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_152_io_a0 = Swapper_120_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_152_io_a1 = Swapper_122_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_153_io_a0 = Swapper_121_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_153_io_a1 = Swapper_123_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_154_io_a0 = Swapper_120_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_154_io_a1 = Swapper_122_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_155_io_a0 = Swapper_121_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_155_io_a1 = Swapper_123_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_156_io_a0 = Swapper_126_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_156_io_a1 = Swapper_124_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_157_io_a0 = Swapper_127_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_157_io_a1 = Swapper_125_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_158_io_a0 = Swapper_126_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_158_io_a1 = Swapper_124_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_159_io_a0 = Swapper_127_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_159_io_a1 = Swapper_125_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_160_io_a0 = Swapper_128_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_160_io_a1 = Swapper_129_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_161_io_a0 = Swapper_128_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_161_io_a1 = Swapper_129_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_162_io_a0 = Swapper_130_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_162_io_a1 = Swapper_131_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_163_io_a0 = Swapper_130_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_163_io_a1 = Swapper_131_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_164_io_a0 = Swapper_133_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_164_io_a1 = Swapper_132_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_165_io_a0 = Swapper_133_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_165_io_a1 = Swapper_132_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_166_io_a0 = Swapper_135_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_166_io_a1 = Swapper_134_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_167_io_a0 = Swapper_135_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_167_io_a1 = Swapper_134_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_168_io_a0 = Swapper_136_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_168_io_a1 = Swapper_137_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_169_io_a0 = Swapper_136_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_169_io_a1 = Swapper_137_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_170_io_a0 = Swapper_138_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_170_io_a1 = Swapper_139_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_171_io_a0 = Swapper_138_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_171_io_a1 = Swapper_139_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_172_io_a0 = Swapper_141_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_172_io_a1 = Swapper_140_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_173_io_a0 = Swapper_141_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_173_io_a1 = Swapper_140_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_174_io_a0 = Swapper_143_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_174_io_a1 = Swapper_142_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_175_io_a0 = Swapper_143_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_175_io_a1 = Swapper_142_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_176_io_a0 = Swapper_144_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_176_io_a1 = Swapper_145_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_177_io_a0 = Swapper_144_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_177_io_a1 = Swapper_145_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_178_io_a0 = Swapper_146_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_178_io_a1 = Swapper_147_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_179_io_a0 = Swapper_146_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_179_io_a1 = Swapper_147_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_180_io_a0 = Swapper_149_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_180_io_a1 = Swapper_148_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_181_io_a0 = Swapper_149_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_181_io_a1 = Swapper_148_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_182_io_a0 = Swapper_151_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_182_io_a1 = Swapper_150_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_183_io_a0 = Swapper_151_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_183_io_a1 = Swapper_150_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_184_io_a0 = Swapper_152_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_184_io_a1 = Swapper_153_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_185_io_a0 = Swapper_152_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_185_io_a1 = Swapper_153_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_186_io_a0 = Swapper_154_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_186_io_a1 = Swapper_155_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_187_io_a0 = Swapper_154_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_187_io_a1 = Swapper_155_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_188_io_a0 = Swapper_157_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_188_io_a1 = Swapper_156_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_189_io_a0 = Swapper_157_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_189_io_a1 = Swapper_156_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_190_io_a0 = Swapper_159_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_190_io_a1 = Swapper_158_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_191_io_a0 = Swapper_159_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_191_io_a1 = Swapper_158_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_192_io_a0 = Swapper_160_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_192_io_a1 = Swapper_164_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_193_io_a0 = Swapper_160_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_193_io_a1 = Swapper_164_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_194_io_a0 = Swapper_161_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_194_io_a1 = Swapper_165_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_195_io_a0 = Swapper_161_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_195_io_a1 = Swapper_165_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_196_io_a0 = Swapper_162_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_196_io_a1 = Swapper_166_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_197_io_a0 = Swapper_162_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_197_io_a1 = Swapper_166_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_198_io_a0 = Swapper_163_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_198_io_a1 = Swapper_167_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_199_io_a0 = Swapper_163_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_199_io_a1 = Swapper_167_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_200_io_a0 = Swapper_172_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_200_io_a1 = Swapper_168_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_201_io_a0 = Swapper_172_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_201_io_a1 = Swapper_168_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_202_io_a0 = Swapper_173_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_202_io_a1 = Swapper_169_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_203_io_a0 = Swapper_173_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_203_io_a1 = Swapper_169_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_204_io_a0 = Swapper_174_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_204_io_a1 = Swapper_170_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_205_io_a0 = Swapper_174_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_205_io_a1 = Swapper_170_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_206_io_a0 = Swapper_175_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_206_io_a1 = Swapper_171_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_207_io_a0 = Swapper_175_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_207_io_a1 = Swapper_171_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_208_io_a0 = Swapper_176_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_208_io_a1 = Swapper_180_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_209_io_a0 = Swapper_176_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_209_io_a1 = Swapper_180_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_210_io_a0 = Swapper_177_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_210_io_a1 = Swapper_181_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_211_io_a0 = Swapper_177_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_211_io_a1 = Swapper_181_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_212_io_a0 = Swapper_178_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_212_io_a1 = Swapper_182_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_213_io_a0 = Swapper_178_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_213_io_a1 = Swapper_182_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_214_io_a0 = Swapper_179_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_214_io_a1 = Swapper_183_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_215_io_a0 = Swapper_179_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_215_io_a1 = Swapper_183_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_216_io_a0 = Swapper_188_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_216_io_a1 = Swapper_184_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_217_io_a0 = Swapper_188_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_217_io_a1 = Swapper_184_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_218_io_a0 = Swapper_189_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_218_io_a1 = Swapper_185_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_219_io_a0 = Swapper_189_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_219_io_a1 = Swapper_185_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_220_io_a0 = Swapper_190_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_220_io_a1 = Swapper_186_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_221_io_a0 = Swapper_190_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_221_io_a1 = Swapper_186_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_222_io_a0 = Swapper_191_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_222_io_a1 = Swapper_187_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_223_io_a0 = Swapper_191_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_223_io_a1 = Swapper_187_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_224_io_a0 = Swapper_192_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_224_io_a1 = Swapper_196_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_225_io_a0 = Swapper_193_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_225_io_a1 = Swapper_197_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_226_io_a0 = Swapper_194_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_226_io_a1 = Swapper_198_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_227_io_a0 = Swapper_195_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_227_io_a1 = Swapper_199_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_228_io_a0 = Swapper_192_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_228_io_a1 = Swapper_196_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_229_io_a0 = Swapper_193_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_229_io_a1 = Swapper_197_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_230_io_a0 = Swapper_194_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_230_io_a1 = Swapper_198_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_231_io_a0 = Swapper_195_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_231_io_a1 = Swapper_199_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_232_io_a0 = Swapper_204_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_232_io_a1 = Swapper_200_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_233_io_a0 = Swapper_205_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_233_io_a1 = Swapper_201_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_234_io_a0 = Swapper_206_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_234_io_a1 = Swapper_202_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_235_io_a0 = Swapper_207_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_235_io_a1 = Swapper_203_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_236_io_a0 = Swapper_204_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_236_io_a1 = Swapper_200_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_237_io_a0 = Swapper_205_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_237_io_a1 = Swapper_201_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_238_io_a0 = Swapper_206_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_238_io_a1 = Swapper_202_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_239_io_a0 = Swapper_207_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_239_io_a1 = Swapper_203_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_240_io_a0 = Swapper_208_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_240_io_a1 = Swapper_212_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_241_io_a0 = Swapper_209_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_241_io_a1 = Swapper_213_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_242_io_a0 = Swapper_210_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_242_io_a1 = Swapper_214_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_243_io_a0 = Swapper_211_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_243_io_a1 = Swapper_215_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_244_io_a0 = Swapper_208_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_244_io_a1 = Swapper_212_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_245_io_a0 = Swapper_209_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_245_io_a1 = Swapper_213_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_246_io_a0 = Swapper_210_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_246_io_a1 = Swapper_214_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_247_io_a0 = Swapper_211_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_247_io_a1 = Swapper_215_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_248_io_a0 = Swapper_220_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_248_io_a1 = Swapper_216_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_249_io_a0 = Swapper_221_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_249_io_a1 = Swapper_217_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_250_io_a0 = Swapper_222_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_250_io_a1 = Swapper_218_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_251_io_a0 = Swapper_223_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_251_io_a1 = Swapper_219_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_252_io_a0 = Swapper_220_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_252_io_a1 = Swapper_216_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_253_io_a0 = Swapper_221_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_253_io_a1 = Swapper_217_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_254_io_a0 = Swapper_222_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_254_io_a1 = Swapper_218_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_255_io_a0 = Swapper_223_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_255_io_a1 = Swapper_219_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_256_io_a0 = Swapper_224_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_256_io_a1 = Swapper_226_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_257_io_a0 = Swapper_225_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_257_io_a1 = Swapper_227_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_258_io_a0 = Swapper_224_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_258_io_a1 = Swapper_226_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_259_io_a0 = Swapper_225_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_259_io_a1 = Swapper_227_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_260_io_a0 = Swapper_228_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_260_io_a1 = Swapper_230_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_261_io_a0 = Swapper_229_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_261_io_a1 = Swapper_231_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_262_io_a0 = Swapper_228_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_262_io_a1 = Swapper_230_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_263_io_a0 = Swapper_229_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_263_io_a1 = Swapper_231_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_264_io_a0 = Swapper_234_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_264_io_a1 = Swapper_232_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_265_io_a0 = Swapper_235_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_265_io_a1 = Swapper_233_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_266_io_a0 = Swapper_234_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_266_io_a1 = Swapper_232_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_267_io_a0 = Swapper_235_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_267_io_a1 = Swapper_233_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_268_io_a0 = Swapper_238_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_268_io_a1 = Swapper_236_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_269_io_a0 = Swapper_239_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_269_io_a1 = Swapper_237_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_270_io_a0 = Swapper_238_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_270_io_a1 = Swapper_236_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_271_io_a0 = Swapper_239_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_271_io_a1 = Swapper_237_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_272_io_a0 = Swapper_240_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_272_io_a1 = Swapper_242_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_273_io_a0 = Swapper_241_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_273_io_a1 = Swapper_243_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_274_io_a0 = Swapper_240_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_274_io_a1 = Swapper_242_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_275_io_a0 = Swapper_241_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_275_io_a1 = Swapper_243_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_276_io_a0 = Swapper_244_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_276_io_a1 = Swapper_246_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_277_io_a0 = Swapper_245_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_277_io_a1 = Swapper_247_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_278_io_a0 = Swapper_244_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_278_io_a1 = Swapper_246_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_279_io_a0 = Swapper_245_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_279_io_a1 = Swapper_247_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_280_io_a0 = Swapper_250_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_280_io_a1 = Swapper_248_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_281_io_a0 = Swapper_251_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_281_io_a1 = Swapper_249_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_282_io_a0 = Swapper_250_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_282_io_a1 = Swapper_248_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_283_io_a0 = Swapper_251_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_283_io_a1 = Swapper_249_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_284_io_a0 = Swapper_254_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_284_io_a1 = Swapper_252_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_285_io_a0 = Swapper_255_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_285_io_a1 = Swapper_253_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_286_io_a0 = Swapper_254_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_286_io_a1 = Swapper_252_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_287_io_a0 = Swapper_255_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_287_io_a1 = Swapper_253_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_288_io_a0 = Swapper_256_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_288_io_a1 = Swapper_257_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_289_io_a0 = Swapper_256_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_289_io_a1 = Swapper_257_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_290_io_a0 = Swapper_258_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_290_io_a1 = Swapper_259_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_291_io_a0 = Swapper_258_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_291_io_a1 = Swapper_259_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_292_io_a0 = Swapper_260_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_292_io_a1 = Swapper_261_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_293_io_a0 = Swapper_260_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_293_io_a1 = Swapper_261_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_294_io_a0 = Swapper_262_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_294_io_a1 = Swapper_263_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_295_io_a0 = Swapper_262_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_295_io_a1 = Swapper_263_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_296_io_a0 = Swapper_265_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_296_io_a1 = Swapper_264_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_297_io_a0 = Swapper_265_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_297_io_a1 = Swapper_264_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_298_io_a0 = Swapper_267_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_298_io_a1 = Swapper_266_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_299_io_a0 = Swapper_267_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_299_io_a1 = Swapper_266_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_300_io_a0 = Swapper_269_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_300_io_a1 = Swapper_268_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_301_io_a0 = Swapper_269_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_301_io_a1 = Swapper_268_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_302_io_a0 = Swapper_271_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_302_io_a1 = Swapper_270_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_303_io_a0 = Swapper_271_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_303_io_a1 = Swapper_270_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_304_io_a0 = Swapper_272_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_304_io_a1 = Swapper_273_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_305_io_a0 = Swapper_272_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_305_io_a1 = Swapper_273_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_306_io_a0 = Swapper_274_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_306_io_a1 = Swapper_275_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_307_io_a0 = Swapper_274_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_307_io_a1 = Swapper_275_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_308_io_a0 = Swapper_276_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_308_io_a1 = Swapper_277_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_309_io_a0 = Swapper_276_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_309_io_a1 = Swapper_277_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_310_io_a0 = Swapper_278_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_310_io_a1 = Swapper_279_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_311_io_a0 = Swapper_278_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_311_io_a1 = Swapper_279_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_312_io_a0 = Swapper_281_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_312_io_a1 = Swapper_280_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_313_io_a0 = Swapper_281_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_313_io_a1 = Swapper_280_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_314_io_a0 = Swapper_283_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_314_io_a1 = Swapper_282_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_315_io_a0 = Swapper_283_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_315_io_a1 = Swapper_282_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_316_io_a0 = Swapper_285_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_316_io_a1 = Swapper_284_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_317_io_a0 = Swapper_285_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_317_io_a1 = Swapper_284_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_318_io_a0 = Swapper_287_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_318_io_a1 = Swapper_286_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_319_io_a0 = Swapper_287_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_319_io_a1 = Swapper_286_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_320_io_a0 = Swapper_288_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_320_io_a1 = Swapper_296_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_321_io_a0 = Swapper_288_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_321_io_a1 = Swapper_296_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_322_io_a0 = Swapper_289_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_322_io_a1 = Swapper_297_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_323_io_a0 = Swapper_289_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_323_io_a1 = Swapper_297_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_324_io_a0 = Swapper_290_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_324_io_a1 = Swapper_298_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_325_io_a0 = Swapper_290_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_325_io_a1 = Swapper_298_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_326_io_a0 = Swapper_291_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_326_io_a1 = Swapper_299_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_327_io_a0 = Swapper_291_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_327_io_a1 = Swapper_299_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_328_io_a0 = Swapper_292_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_328_io_a1 = Swapper_300_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_329_io_a0 = Swapper_292_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_329_io_a1 = Swapper_300_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_330_io_a0 = Swapper_293_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_330_io_a1 = Swapper_301_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_331_io_a0 = Swapper_293_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_331_io_a1 = Swapper_301_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_332_io_a0 = Swapper_294_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_332_io_a1 = Swapper_302_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_333_io_a0 = Swapper_294_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_333_io_a1 = Swapper_302_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_334_io_a0 = Swapper_295_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_334_io_a1 = Swapper_303_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_335_io_a0 = Swapper_295_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_335_io_a1 = Swapper_303_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_336_io_a0 = Swapper_312_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_336_io_a1 = Swapper_304_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_337_io_a0 = Swapper_312_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_337_io_a1 = Swapper_304_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_338_io_a0 = Swapper_313_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_338_io_a1 = Swapper_305_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_339_io_a0 = Swapper_313_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_339_io_a1 = Swapper_305_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_340_io_a0 = Swapper_314_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_340_io_a1 = Swapper_306_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_341_io_a0 = Swapper_314_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_341_io_a1 = Swapper_306_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_342_io_a0 = Swapper_315_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_342_io_a1 = Swapper_307_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_343_io_a0 = Swapper_315_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_343_io_a1 = Swapper_307_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_344_io_a0 = Swapper_316_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_344_io_a1 = Swapper_308_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_345_io_a0 = Swapper_316_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_345_io_a1 = Swapper_308_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_346_io_a0 = Swapper_317_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_346_io_a1 = Swapper_309_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_347_io_a0 = Swapper_317_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_347_io_a1 = Swapper_309_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_348_io_a0 = Swapper_318_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_348_io_a1 = Swapper_310_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_349_io_a0 = Swapper_318_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_349_io_a1 = Swapper_310_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_350_io_a0 = Swapper_319_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_350_io_a1 = Swapper_311_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_351_io_a0 = Swapper_319_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_351_io_a1 = Swapper_311_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_352_io_a0 = Swapper_320_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_352_io_a1 = Swapper_328_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_353_io_a0 = Swapper_321_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_353_io_a1 = Swapper_329_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_354_io_a0 = Swapper_322_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_354_io_a1 = Swapper_330_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_355_io_a0 = Swapper_323_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_355_io_a1 = Swapper_331_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_356_io_a0 = Swapper_324_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_356_io_a1 = Swapper_332_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_357_io_a0 = Swapper_325_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_357_io_a1 = Swapper_333_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_358_io_a0 = Swapper_326_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_358_io_a1 = Swapper_334_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_359_io_a0 = Swapper_327_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_359_io_a1 = Swapper_335_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_360_io_a0 = Swapper_320_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_360_io_a1 = Swapper_328_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_361_io_a0 = Swapper_321_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_361_io_a1 = Swapper_329_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_362_io_a0 = Swapper_322_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_362_io_a1 = Swapper_330_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_363_io_a0 = Swapper_323_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_363_io_a1 = Swapper_331_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_364_io_a0 = Swapper_324_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_364_io_a1 = Swapper_332_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_365_io_a0 = Swapper_325_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_365_io_a1 = Swapper_333_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_366_io_a0 = Swapper_326_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_366_io_a1 = Swapper_334_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_367_io_a0 = Swapper_327_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_367_io_a1 = Swapper_335_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_368_io_a0 = Swapper_344_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_368_io_a1 = Swapper_336_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_369_io_a0 = Swapper_345_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_369_io_a1 = Swapper_337_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_370_io_a0 = Swapper_346_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_370_io_a1 = Swapper_338_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_371_io_a0 = Swapper_347_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_371_io_a1 = Swapper_339_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_372_io_a0 = Swapper_348_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_372_io_a1 = Swapper_340_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_373_io_a0 = Swapper_349_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_373_io_a1 = Swapper_341_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_374_io_a0 = Swapper_350_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_374_io_a1 = Swapper_342_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_375_io_a0 = Swapper_351_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_375_io_a1 = Swapper_343_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_376_io_a0 = Swapper_344_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_376_io_a1 = Swapper_336_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_377_io_a0 = Swapper_345_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_377_io_a1 = Swapper_337_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_378_io_a0 = Swapper_346_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_378_io_a1 = Swapper_338_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_379_io_a0 = Swapper_347_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_379_io_a1 = Swapper_339_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_380_io_a0 = Swapper_348_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_380_io_a1 = Swapper_340_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_381_io_a0 = Swapper_349_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_381_io_a1 = Swapper_341_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_382_io_a0 = Swapper_350_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_382_io_a1 = Swapper_342_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_383_io_a0 = Swapper_351_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_383_io_a1 = Swapper_343_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_384_io_a0 = Swapper_352_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_384_io_a1 = Swapper_356_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_385_io_a0 = Swapper_353_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_385_io_a1 = Swapper_357_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_386_io_a0 = Swapper_354_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_386_io_a1 = Swapper_358_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_387_io_a0 = Swapper_355_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_387_io_a1 = Swapper_359_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_388_io_a0 = Swapper_352_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_388_io_a1 = Swapper_356_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_389_io_a0 = Swapper_353_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_389_io_a1 = Swapper_357_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_390_io_a0 = Swapper_354_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_390_io_a1 = Swapper_358_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_391_io_a0 = Swapper_355_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_391_io_a1 = Swapper_359_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_392_io_a0 = Swapper_360_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_392_io_a1 = Swapper_364_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_393_io_a0 = Swapper_361_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_393_io_a1 = Swapper_365_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_394_io_a0 = Swapper_362_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_394_io_a1 = Swapper_366_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_395_io_a0 = Swapper_363_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_395_io_a1 = Swapper_367_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_396_io_a0 = Swapper_360_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_396_io_a1 = Swapper_364_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_397_io_a0 = Swapper_361_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_397_io_a1 = Swapper_365_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_398_io_a0 = Swapper_362_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_398_io_a1 = Swapper_366_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_399_io_a0 = Swapper_363_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_399_io_a1 = Swapper_367_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_400_io_a0 = Swapper_372_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_400_io_a1 = Swapper_368_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_401_io_a0 = Swapper_373_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_401_io_a1 = Swapper_369_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_402_io_a0 = Swapper_374_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_402_io_a1 = Swapper_370_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_403_io_a0 = Swapper_375_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_403_io_a1 = Swapper_371_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_404_io_a0 = Swapper_372_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_404_io_a1 = Swapper_368_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_405_io_a0 = Swapper_373_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_405_io_a1 = Swapper_369_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_406_io_a0 = Swapper_374_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_406_io_a1 = Swapper_370_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_407_io_a0 = Swapper_375_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_407_io_a1 = Swapper_371_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_408_io_a0 = Swapper_380_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_408_io_a1 = Swapper_376_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_409_io_a0 = Swapper_381_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_409_io_a1 = Swapper_377_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_410_io_a0 = Swapper_382_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_410_io_a1 = Swapper_378_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_411_io_a0 = Swapper_383_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_411_io_a1 = Swapper_379_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_412_io_a0 = Swapper_380_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_412_io_a1 = Swapper_376_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_413_io_a0 = Swapper_381_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_413_io_a1 = Swapper_377_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_414_io_a0 = Swapper_382_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_414_io_a1 = Swapper_378_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_415_io_a0 = Swapper_383_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_415_io_a1 = Swapper_379_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_416_io_a0 = Swapper_384_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_416_io_a1 = Swapper_386_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_417_io_a0 = Swapper_385_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_417_io_a1 = Swapper_387_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_418_io_a0 = Swapper_384_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_418_io_a1 = Swapper_386_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_419_io_a0 = Swapper_385_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_419_io_a1 = Swapper_387_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_420_io_a0 = Swapper_388_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_420_io_a1 = Swapper_390_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_421_io_a0 = Swapper_389_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_421_io_a1 = Swapper_391_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_422_io_a0 = Swapper_388_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_422_io_a1 = Swapper_390_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_423_io_a0 = Swapper_389_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_423_io_a1 = Swapper_391_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_424_io_a0 = Swapper_392_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_424_io_a1 = Swapper_394_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_425_io_a0 = Swapper_393_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_425_io_a1 = Swapper_395_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_426_io_a0 = Swapper_392_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_426_io_a1 = Swapper_394_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_427_io_a0 = Swapper_393_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_427_io_a1 = Swapper_395_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_428_io_a0 = Swapper_396_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_428_io_a1 = Swapper_398_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_429_io_a0 = Swapper_397_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_429_io_a1 = Swapper_399_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_430_io_a0 = Swapper_396_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_430_io_a1 = Swapper_398_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_431_io_a0 = Swapper_397_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_431_io_a1 = Swapper_399_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_432_io_a0 = Swapper_402_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_432_io_a1 = Swapper_400_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_433_io_a0 = Swapper_403_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_433_io_a1 = Swapper_401_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_434_io_a0 = Swapper_402_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_434_io_a1 = Swapper_400_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_435_io_a0 = Swapper_403_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_435_io_a1 = Swapper_401_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_436_io_a0 = Swapper_406_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_436_io_a1 = Swapper_404_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_437_io_a0 = Swapper_407_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_437_io_a1 = Swapper_405_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_438_io_a0 = Swapper_406_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_438_io_a1 = Swapper_404_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_439_io_a0 = Swapper_407_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_439_io_a1 = Swapper_405_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_440_io_a0 = Swapper_410_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_440_io_a1 = Swapper_408_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_441_io_a0 = Swapper_411_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_441_io_a1 = Swapper_409_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_442_io_a0 = Swapper_410_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_442_io_a1 = Swapper_408_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_443_io_a0 = Swapper_411_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_443_io_a1 = Swapper_409_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_444_io_a0 = Swapper_414_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_444_io_a1 = Swapper_412_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_445_io_a0 = Swapper_415_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_445_io_a1 = Swapper_413_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_446_io_a0 = Swapper_414_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_446_io_a1 = Swapper_412_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_447_io_a0 = Swapper_415_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_447_io_a1 = Swapper_413_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_448_io_a0 = Swapper_416_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_448_io_a1 = Swapper_417_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_449_io_a0 = Swapper_416_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_449_io_a1 = Swapper_417_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_450_io_a0 = Swapper_418_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_450_io_a1 = Swapper_419_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_451_io_a0 = Swapper_418_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_451_io_a1 = Swapper_419_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_452_io_a0 = Swapper_420_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_452_io_a1 = Swapper_421_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_453_io_a0 = Swapper_420_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_453_io_a1 = Swapper_421_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_454_io_a0 = Swapper_422_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_454_io_a1 = Swapper_423_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_455_io_a0 = Swapper_422_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_455_io_a1 = Swapper_423_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_456_io_a0 = Swapper_424_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_456_io_a1 = Swapper_425_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_457_io_a0 = Swapper_424_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_457_io_a1 = Swapper_425_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_458_io_a0 = Swapper_426_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_458_io_a1 = Swapper_427_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_459_io_a0 = Swapper_426_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_459_io_a1 = Swapper_427_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_460_io_a0 = Swapper_428_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_460_io_a1 = Swapper_429_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_461_io_a0 = Swapper_428_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_461_io_a1 = Swapper_429_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_462_io_a0 = Swapper_430_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_462_io_a1 = Swapper_431_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_463_io_a0 = Swapper_430_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_463_io_a1 = Swapper_431_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_464_io_a0 = Swapper_433_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_464_io_a1 = Swapper_432_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_465_io_a0 = Swapper_433_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_465_io_a1 = Swapper_432_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_466_io_a0 = Swapper_435_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_466_io_a1 = Swapper_434_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_467_io_a0 = Swapper_435_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_467_io_a1 = Swapper_434_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_468_io_a0 = Swapper_437_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_468_io_a1 = Swapper_436_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_469_io_a0 = Swapper_437_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_469_io_a1 = Swapper_436_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_470_io_a0 = Swapper_439_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_470_io_a1 = Swapper_438_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_471_io_a0 = Swapper_439_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_471_io_a1 = Swapper_438_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_472_io_a0 = Swapper_441_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_472_io_a1 = Swapper_440_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_473_io_a0 = Swapper_441_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_473_io_a1 = Swapper_440_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_474_io_a0 = Swapper_443_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_474_io_a1 = Swapper_442_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_475_io_a0 = Swapper_443_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_475_io_a1 = Swapper_442_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_476_io_a0 = Swapper_445_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_476_io_a1 = Swapper_444_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_477_io_a0 = Swapper_445_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_477_io_a1 = Swapper_444_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_478_io_a0 = Swapper_447_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_478_io_a1 = Swapper_446_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_479_io_a0 = Swapper_447_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_479_io_a1 = Swapper_446_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_480_io_a0 = Swapper_448_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_480_io_a1 = Swapper_464_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_481_io_a0 = Swapper_448_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_481_io_a1 = Swapper_464_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_482_io_a0 = Swapper_449_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_482_io_a1 = Swapper_465_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_483_io_a0 = Swapper_449_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_483_io_a1 = Swapper_465_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_484_io_a0 = Swapper_450_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_484_io_a1 = Swapper_466_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_485_io_a0 = Swapper_450_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_485_io_a1 = Swapper_466_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_486_io_a0 = Swapper_451_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_486_io_a1 = Swapper_467_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_487_io_a0 = Swapper_451_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_487_io_a1 = Swapper_467_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_488_io_a0 = Swapper_452_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_488_io_a1 = Swapper_468_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_489_io_a0 = Swapper_452_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_489_io_a1 = Swapper_468_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_490_io_a0 = Swapper_453_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_490_io_a1 = Swapper_469_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_491_io_a0 = Swapper_453_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_491_io_a1 = Swapper_469_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_492_io_a0 = Swapper_454_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_492_io_a1 = Swapper_470_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_493_io_a0 = Swapper_454_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_493_io_a1 = Swapper_470_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_494_io_a0 = Swapper_455_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_494_io_a1 = Swapper_471_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_495_io_a0 = Swapper_455_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_495_io_a1 = Swapper_471_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_496_io_a0 = Swapper_456_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_496_io_a1 = Swapper_472_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_497_io_a0 = Swapper_456_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_497_io_a1 = Swapper_472_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_498_io_a0 = Swapper_457_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_498_io_a1 = Swapper_473_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_499_io_a0 = Swapper_457_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_499_io_a1 = Swapper_473_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_500_io_a0 = Swapper_458_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_500_io_a1 = Swapper_474_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_501_io_a0 = Swapper_458_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_501_io_a1 = Swapper_474_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_502_io_a0 = Swapper_459_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_502_io_a1 = Swapper_475_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_503_io_a0 = Swapper_459_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_503_io_a1 = Swapper_475_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_504_io_a0 = Swapper_460_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_504_io_a1 = Swapper_476_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_505_io_a0 = Swapper_460_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_505_io_a1 = Swapper_476_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_506_io_a0 = Swapper_461_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_506_io_a1 = Swapper_477_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_507_io_a0 = Swapper_461_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_507_io_a1 = Swapper_477_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_508_io_a0 = Swapper_462_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_508_io_a1 = Swapper_478_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_509_io_a0 = Swapper_462_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_509_io_a1 = Swapper_478_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_510_io_a0 = Swapper_463_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_510_io_a1 = Swapper_479_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_511_io_a0 = Swapper_463_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_511_io_a1 = Swapper_479_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_512_io_a0 = Swapper_480_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_512_io_a1 = Swapper_496_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_513_io_a0 = Swapper_481_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_513_io_a1 = Swapper_497_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_514_io_a0 = Swapper_482_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_514_io_a1 = Swapper_498_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_515_io_a0 = Swapper_483_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_515_io_a1 = Swapper_499_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_516_io_a0 = Swapper_484_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_516_io_a1 = Swapper_500_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_517_io_a0 = Swapper_485_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_517_io_a1 = Swapper_501_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_518_io_a0 = Swapper_486_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_518_io_a1 = Swapper_502_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_519_io_a0 = Swapper_487_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_519_io_a1 = Swapper_503_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_520_io_a0 = Swapper_488_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_520_io_a1 = Swapper_504_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_521_io_a0 = Swapper_489_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_521_io_a1 = Swapper_505_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_522_io_a0 = Swapper_490_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_522_io_a1 = Swapper_506_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_523_io_a0 = Swapper_491_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_523_io_a1 = Swapper_507_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_524_io_a0 = Swapper_492_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_524_io_a1 = Swapper_508_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_525_io_a0 = Swapper_493_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_525_io_a1 = Swapper_509_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_526_io_a0 = Swapper_494_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_526_io_a1 = Swapper_510_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_527_io_a0 = Swapper_495_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_527_io_a1 = Swapper_511_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_528_io_a0 = Swapper_480_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_528_io_a1 = Swapper_496_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_529_io_a0 = Swapper_481_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_529_io_a1 = Swapper_497_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_530_io_a0 = Swapper_482_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_530_io_a1 = Swapper_498_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_531_io_a0 = Swapper_483_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_531_io_a1 = Swapper_499_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_532_io_a0 = Swapper_484_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_532_io_a1 = Swapper_500_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_533_io_a0 = Swapper_485_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_533_io_a1 = Swapper_501_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_534_io_a0 = Swapper_486_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_534_io_a1 = Swapper_502_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_535_io_a0 = Swapper_487_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_535_io_a1 = Swapper_503_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_536_io_a0 = Swapper_488_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_536_io_a1 = Swapper_504_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_537_io_a0 = Swapper_489_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_537_io_a1 = Swapper_505_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_538_io_a0 = Swapper_490_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_538_io_a1 = Swapper_506_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_539_io_a0 = Swapper_491_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_539_io_a1 = Swapper_507_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_540_io_a0 = Swapper_492_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_540_io_a1 = Swapper_508_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_541_io_a0 = Swapper_493_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_541_io_a1 = Swapper_509_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_542_io_a0 = Swapper_494_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_542_io_a1 = Swapper_510_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_543_io_a0 = Swapper_495_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_543_io_a1 = Swapper_511_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_544_io_a0 = Swapper_512_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_544_io_a1 = Swapper_520_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_545_io_a0 = Swapper_513_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_545_io_a1 = Swapper_521_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_546_io_a0 = Swapper_514_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_546_io_a1 = Swapper_522_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_547_io_a0 = Swapper_515_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_547_io_a1 = Swapper_523_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_548_io_a0 = Swapper_516_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_548_io_a1 = Swapper_524_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_549_io_a0 = Swapper_517_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_549_io_a1 = Swapper_525_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_550_io_a0 = Swapper_518_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_550_io_a1 = Swapper_526_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_551_io_a0 = Swapper_519_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_551_io_a1 = Swapper_527_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_552_io_a0 = Swapper_512_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_552_io_a1 = Swapper_520_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_553_io_a0 = Swapper_513_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_553_io_a1 = Swapper_521_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_554_io_a0 = Swapper_514_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_554_io_a1 = Swapper_522_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_555_io_a0 = Swapper_515_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_555_io_a1 = Swapper_523_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_556_io_a0 = Swapper_516_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_556_io_a1 = Swapper_524_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_557_io_a0 = Swapper_517_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_557_io_a1 = Swapper_525_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_558_io_a0 = Swapper_518_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_558_io_a1 = Swapper_526_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_559_io_a0 = Swapper_519_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_559_io_a1 = Swapper_527_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_560_io_a0 = Swapper_528_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_560_io_a1 = Swapper_536_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_561_io_a0 = Swapper_529_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_561_io_a1 = Swapper_537_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_562_io_a0 = Swapper_530_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_562_io_a1 = Swapper_538_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_563_io_a0 = Swapper_531_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_563_io_a1 = Swapper_539_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_564_io_a0 = Swapper_532_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_564_io_a1 = Swapper_540_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_565_io_a0 = Swapper_533_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_565_io_a1 = Swapper_541_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_566_io_a0 = Swapper_534_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_566_io_a1 = Swapper_542_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_567_io_a0 = Swapper_535_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_567_io_a1 = Swapper_543_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_568_io_a0 = Swapper_528_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_568_io_a1 = Swapper_536_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_569_io_a0 = Swapper_529_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_569_io_a1 = Swapper_537_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_570_io_a0 = Swapper_530_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_570_io_a1 = Swapper_538_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_571_io_a0 = Swapper_531_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_571_io_a1 = Swapper_539_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_572_io_a0 = Swapper_532_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_572_io_a1 = Swapper_540_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_573_io_a0 = Swapper_533_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_573_io_a1 = Swapper_541_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_574_io_a0 = Swapper_534_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_574_io_a1 = Swapper_542_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_575_io_a0 = Swapper_535_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_575_io_a1 = Swapper_543_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_576_io_a0 = Swapper_544_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_576_io_a1 = Swapper_548_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_577_io_a0 = Swapper_545_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_577_io_a1 = Swapper_549_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_578_io_a0 = Swapper_546_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_578_io_a1 = Swapper_550_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_579_io_a0 = Swapper_547_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_579_io_a1 = Swapper_551_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_580_io_a0 = Swapper_544_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_580_io_a1 = Swapper_548_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_581_io_a0 = Swapper_545_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_581_io_a1 = Swapper_549_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_582_io_a0 = Swapper_546_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_582_io_a1 = Swapper_550_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_583_io_a0 = Swapper_547_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_583_io_a1 = Swapper_551_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_584_io_a0 = Swapper_552_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_584_io_a1 = Swapper_556_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_585_io_a0 = Swapper_553_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_585_io_a1 = Swapper_557_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_586_io_a0 = Swapper_554_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_586_io_a1 = Swapper_558_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_587_io_a0 = Swapper_555_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_587_io_a1 = Swapper_559_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_588_io_a0 = Swapper_552_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_588_io_a1 = Swapper_556_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_589_io_a0 = Swapper_553_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_589_io_a1 = Swapper_557_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_590_io_a0 = Swapper_554_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_590_io_a1 = Swapper_558_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_591_io_a0 = Swapper_555_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_591_io_a1 = Swapper_559_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_592_io_a0 = Swapper_560_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_592_io_a1 = Swapper_564_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_593_io_a0 = Swapper_561_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_593_io_a1 = Swapper_565_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_594_io_a0 = Swapper_562_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_594_io_a1 = Swapper_566_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_595_io_a0 = Swapper_563_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_595_io_a1 = Swapper_567_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_596_io_a0 = Swapper_560_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_596_io_a1 = Swapper_564_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_597_io_a0 = Swapper_561_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_597_io_a1 = Swapper_565_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_598_io_a0 = Swapper_562_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_598_io_a1 = Swapper_566_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_599_io_a0 = Swapper_563_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_599_io_a1 = Swapper_567_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_600_io_a0 = Swapper_568_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_600_io_a1 = Swapper_572_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_601_io_a0 = Swapper_569_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_601_io_a1 = Swapper_573_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_602_io_a0 = Swapper_570_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_602_io_a1 = Swapper_574_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_603_io_a0 = Swapper_571_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_603_io_a1 = Swapper_575_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_604_io_a0 = Swapper_568_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_604_io_a1 = Swapper_572_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_605_io_a0 = Swapper_569_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_605_io_a1 = Swapper_573_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_606_io_a0 = Swapper_570_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_606_io_a1 = Swapper_574_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_607_io_a0 = Swapper_571_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_607_io_a1 = Swapper_575_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_608_io_a0 = Swapper_576_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_608_io_a1 = Swapper_578_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_609_io_a0 = Swapper_577_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_609_io_a1 = Swapper_579_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_610_io_a0 = Swapper_576_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_610_io_a1 = Swapper_578_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_611_io_a0 = Swapper_577_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_611_io_a1 = Swapper_579_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_612_io_a0 = Swapper_580_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_612_io_a1 = Swapper_582_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_613_io_a0 = Swapper_581_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_613_io_a1 = Swapper_583_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_614_io_a0 = Swapper_580_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_614_io_a1 = Swapper_582_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_615_io_a0 = Swapper_581_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_615_io_a1 = Swapper_583_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_616_io_a0 = Swapper_584_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_616_io_a1 = Swapper_586_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_617_io_a0 = Swapper_585_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_617_io_a1 = Swapper_587_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_618_io_a0 = Swapper_584_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_618_io_a1 = Swapper_586_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_619_io_a0 = Swapper_585_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_619_io_a1 = Swapper_587_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_620_io_a0 = Swapper_588_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_620_io_a1 = Swapper_590_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_621_io_a0 = Swapper_589_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_621_io_a1 = Swapper_591_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_622_io_a0 = Swapper_588_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_622_io_a1 = Swapper_590_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_623_io_a0 = Swapper_589_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_623_io_a1 = Swapper_591_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_624_io_a0 = Swapper_592_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_624_io_a1 = Swapper_594_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_625_io_a0 = Swapper_593_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_625_io_a1 = Swapper_595_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_626_io_a0 = Swapper_592_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_626_io_a1 = Swapper_594_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_627_io_a0 = Swapper_593_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_627_io_a1 = Swapper_595_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_628_io_a0 = Swapper_596_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_628_io_a1 = Swapper_598_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_629_io_a0 = Swapper_597_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_629_io_a1 = Swapper_599_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_630_io_a0 = Swapper_596_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_630_io_a1 = Swapper_598_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_631_io_a0 = Swapper_597_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_631_io_a1 = Swapper_599_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_632_io_a0 = Swapper_600_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_632_io_a1 = Swapper_602_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_633_io_a0 = Swapper_601_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_633_io_a1 = Swapper_603_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_634_io_a0 = Swapper_600_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_634_io_a1 = Swapper_602_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_635_io_a0 = Swapper_601_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_635_io_a1 = Swapper_603_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_636_io_a0 = Swapper_604_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_636_io_a1 = Swapper_606_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_637_io_a0 = Swapper_605_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_637_io_a1 = Swapper_607_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_638_io_a0 = Swapper_604_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_638_io_a1 = Swapper_606_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_639_io_a0 = Swapper_605_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_639_io_a1 = Swapper_607_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_640_io_a0 = Swapper_608_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_640_io_a1 = Swapper_609_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_641_io_a0 = Swapper_608_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_641_io_a1 = Swapper_609_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_642_io_a0 = Swapper_610_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_642_io_a1 = Swapper_611_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_643_io_a0 = Swapper_610_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_643_io_a1 = Swapper_611_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_644_io_a0 = Swapper_612_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_644_io_a1 = Swapper_613_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_645_io_a0 = Swapper_612_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_645_io_a1 = Swapper_613_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_646_io_a0 = Swapper_614_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_646_io_a1 = Swapper_615_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_647_io_a0 = Swapper_614_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_647_io_a1 = Swapper_615_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_648_io_a0 = Swapper_616_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_648_io_a1 = Swapper_617_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_649_io_a0 = Swapper_616_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_649_io_a1 = Swapper_617_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_650_io_a0 = Swapper_618_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_650_io_a1 = Swapper_619_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_651_io_a0 = Swapper_618_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_651_io_a1 = Swapper_619_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_652_io_a0 = Swapper_620_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_652_io_a1 = Swapper_621_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_653_io_a0 = Swapper_620_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_653_io_a1 = Swapper_621_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_654_io_a0 = Swapper_622_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_654_io_a1 = Swapper_623_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_655_io_a0 = Swapper_622_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_655_io_a1 = Swapper_623_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_656_io_a0 = Swapper_624_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_656_io_a1 = Swapper_625_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_657_io_a0 = Swapper_624_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_657_io_a1 = Swapper_625_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_658_io_a0 = Swapper_626_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_658_io_a1 = Swapper_627_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_659_io_a0 = Swapper_626_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_659_io_a1 = Swapper_627_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_660_io_a0 = Swapper_628_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_660_io_a1 = Swapper_629_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_661_io_a0 = Swapper_628_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_661_io_a1 = Swapper_629_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_662_io_a0 = Swapper_630_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_662_io_a1 = Swapper_631_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_663_io_a0 = Swapper_630_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_663_io_a1 = Swapper_631_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_664_io_a0 = Swapper_632_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_664_io_a1 = Swapper_633_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_665_io_a0 = Swapper_632_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_665_io_a1 = Swapper_633_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_666_io_a0 = Swapper_634_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_666_io_a1 = Swapper_635_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_667_io_a0 = Swapper_634_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_667_io_a1 = Swapper_635_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_668_io_a0 = Swapper_636_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_668_io_a1 = Swapper_637_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_669_io_a0 = Swapper_636_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_669_io_a1 = Swapper_637_io_z1; // @[bitonic_sort.scala 33:19]
  assign Swapper_670_io_a0 = Swapper_638_io_z0; // @[bitonic_sort.scala 32:19]
  assign Swapper_670_io_a1 = Swapper_639_io_z0; // @[bitonic_sort.scala 33:19]
  assign Swapper_671_io_a0 = Swapper_638_io_z1; // @[bitonic_sort.scala 32:19]
  assign Swapper_671_io_a1 = Swapper_639_io_z1; // @[bitonic_sort.scala 33:19]

initial begin
   $vcdplusfile("/nfs/site/disks/scl.work.37/ppt/users/smburns/cocotb-pg/agile-hardware-using-verilog/bitonic/tests/foo.vpd");
   $vcdpluson(0);
end
   

endmodule
