module Splitter(
  output        io_mi_ready,
  input         io_mi_valid,
  input  [15:0] io_mi_bits_0,
  input  [15:0] io_mi_bits_1,
  input  [15:0] io_mi_bits_2,
  input  [15:0] io_mi_bits_3,
  input  [15:0] io_mi_bits_4,
  input  [15:0] io_mi_bits_5,
  input  [15:0] io_mi_bits_6,
  input  [15:0] io_mi_bits_7,
  input         io_mi0_ready,
  output        io_mi0_valid,
  output [15:0] io_mi0_bits_0,
  output [15:0] io_mi0_bits_1,
  output [15:0] io_mi0_bits_2,
  output [15:0] io_mi0_bits_3,
  output [15:0] io_mi0_bits_4,
  output [15:0] io_mi0_bits_5,
  output [15:0] io_mi0_bits_6,
  output [15:0] io_mi0_bits_7,
  input         io_mi1_ready,
  output        io_mi1_valid,
  output [15:0] io_mi1_bits_0,
  output [15:0] io_mi1_bits_1,
  output [15:0] io_mi1_bits_2,
  output [15:0] io_mi1_bits_3,
  output [15:0] io_mi1_bits_4,
  output [15:0] io_mi1_bits_5,
  output [15:0] io_mi1_bits_6,
  output [15:0] io_mi1_bits_7
);
  wire  _T; // @[Splitter.scala 19:22]
  assign _T = io_mi_valid & io_mi0_ready; // @[Splitter.scala 19:22]
  assign io_mi_ready = _T & io_mi1_ready; // @[Decoupled.scala 69:20 Splitter.scala 20:17]
  assign io_mi0_valid = _T & io_mi1_ready; // @[Decoupled.scala 53:20 Splitter.scala 21:18]
  assign io_mi0_bits_0 = io_mi_bits_0; // @[Splitter.scala 23:17]
  assign io_mi0_bits_1 = io_mi_bits_1; // @[Splitter.scala 23:17]
  assign io_mi0_bits_2 = io_mi_bits_2; // @[Splitter.scala 23:17]
  assign io_mi0_bits_3 = io_mi_bits_3; // @[Splitter.scala 23:17]
  assign io_mi0_bits_4 = io_mi_bits_4; // @[Splitter.scala 23:17]
  assign io_mi0_bits_5 = io_mi_bits_5; // @[Splitter.scala 23:17]
  assign io_mi0_bits_6 = io_mi_bits_6; // @[Splitter.scala 23:17]
  assign io_mi0_bits_7 = io_mi_bits_7; // @[Splitter.scala 23:17]
  assign io_mi1_valid = _T & io_mi1_ready; // @[Decoupled.scala 53:20 Splitter.scala 22:18]
  assign io_mi1_bits_0 = io_mi_bits_0; // @[Splitter.scala 24:17]
  assign io_mi1_bits_1 = io_mi_bits_1; // @[Splitter.scala 24:17]
  assign io_mi1_bits_2 = io_mi_bits_2; // @[Splitter.scala 24:17]
  assign io_mi1_bits_3 = io_mi_bits_3; // @[Splitter.scala 24:17]
  assign io_mi1_bits_4 = io_mi_bits_4; // @[Splitter.scala 24:17]
  assign io_mi1_bits_5 = io_mi_bits_5; // @[Splitter.scala 24:17]
  assign io_mi1_bits_6 = io_mi_bits_6; // @[Splitter.scala 24:17]
  assign io_mi1_bits_7 = io_mi_bits_7; // @[Splitter.scala 24:17]
endmodule
module Frontend(
  input         clock,
  input         reset,
  input         io_start,
  output        io_gi_ready,
  input         io_gi_valid,
  input  [15:0] io_gi_bits_0,
  input  [15:0] io_gi_bits_1,
  input  [15:0] io_gi_bits_2,
  input  [15:0] io_gi_bits_3,
  input  [15:0] io_gi_bits_4,
  input  [15:0] io_gi_bits_5,
  input  [15:0] io_gi_bits_6,
  input  [15:0] io_gi_bits_7,
  output        io_wi_ready,
  input         io_wi_valid,
  input  [15:0] io_wi_bits_0,
  input  [15:0] io_wi_bits_1,
  input  [15:0] io_wi_bits_2,
  input  [15:0] io_wi_bits_3,
  input  [15:0] io_wi_bits_4,
  input  [15:0] io_wi_bits_5,
  input  [15:0] io_wi_bits_6,
  input  [15:0] io_wi_bits_7,
  output        io_a0_ready,
  input         io_a0_valid,
  input  [15:0] io_a0_bits_0,
  input  [15:0] io_a0_bits_1,
  input  [15:0] io_a0_bits_2,
  input  [15:0] io_a0_bits_3,
  input  [15:0] io_a0_bits_4,
  input  [15:0] io_a0_bits_5,
  input  [15:0] io_a0_bits_6,
  input  [15:0] io_a0_bits_7,
  output        io_mi1_ready,
  input         io_mi1_valid,
  input  [15:0] io_mi1_bits_0,
  input  [15:0] io_mi1_bits_1,
  input  [15:0] io_mi1_bits_2,
  input  [15:0] io_mi1_bits_3,
  input  [15:0] io_mi1_bits_4,
  input  [15:0] io_mi1_bits_5,
  input  [15:0] io_mi1_bits_6,
  input  [15:0] io_mi1_bits_7,
  output        io_adj_ready,
  input         io_adj_valid,
  input  [15:0] io_adj_bits_0,
  input  [15:0] io_adj_bits_1,
  input  [15:0] io_adj_bits_2,
  input  [15:0] io_adj_bits_3,
  input  [15:0] io_adj_bits_4,
  input  [15:0] io_adj_bits_5,
  input  [15:0] io_adj_bits_6,
  input  [15:0] io_adj_bits_7,
  input         io_off_ready,
  output        io_off_valid,
  output [15:0] io_off_bits_0,
  output [15:0] io_off_bits_1,
  output [15:0] io_off_bits_2,
  output [15:0] io_off_bits_3,
  output [15:0] io_off_bits_4,
  output [15:0] io_off_bits_5,
  output [15:0] io_off_bits_6,
  output [15:0] io_off_bits_7
);
  reg  phase; // @[Frontend.scala 20:22]
  reg [31:0] _RAND_0;
  reg [1:0] jj; // @[Frontend.scala 21:19]
  reg [31:0] _RAND_1;
  reg [1:0] _T; // @[SliceCounter.scala 7:19]
  reg [31:0] _RAND_2;
  reg [4:0] _T_1; // @[SliceCounter.scala 8:19]
  reg [31:0] _RAND_3;
  reg [4:0] _T_2; // @[SliceCounter.scala 9:19]
  reg [31:0] _RAND_4;
  reg  _T_5; // @[SliceCounter.scala 12:24]
  reg [31:0] _RAND_5;
  reg [15:0] gamma_0_0; // @[Frontend.scala 25:18]
  reg [31:0] _RAND_6;
  reg [15:0] gamma_0_1; // @[Frontend.scala 25:18]
  reg [31:0] _RAND_7;
  reg [15:0] gamma_0_2; // @[Frontend.scala 25:18]
  reg [31:0] _RAND_8;
  reg [15:0] gamma_0_3; // @[Frontend.scala 25:18]
  reg [31:0] _RAND_9;
  reg [15:0] gamma_0_4; // @[Frontend.scala 25:18]
  reg [31:0] _RAND_10;
  reg [15:0] gamma_0_5; // @[Frontend.scala 25:18]
  reg [31:0] _RAND_11;
  reg [15:0] gamma_0_6; // @[Frontend.scala 25:18]
  reg [31:0] _RAND_12;
  reg [15:0] gamma_0_7; // @[Frontend.scala 25:18]
  reg [31:0] _RAND_13;
  reg [15:0] gamma_1_0; // @[Frontend.scala 25:18]
  reg [31:0] _RAND_14;
  reg [15:0] gamma_1_1; // @[Frontend.scala 25:18]
  reg [31:0] _RAND_15;
  reg [15:0] gamma_1_2; // @[Frontend.scala 25:18]
  reg [31:0] _RAND_16;
  reg [15:0] gamma_1_3; // @[Frontend.scala 25:18]
  reg [31:0] _RAND_17;
  reg [15:0] gamma_1_4; // @[Frontend.scala 25:18]
  reg [31:0] _RAND_18;
  reg [15:0] gamma_1_5; // @[Frontend.scala 25:18]
  reg [31:0] _RAND_19;
  reg [15:0] gamma_1_6; // @[Frontend.scala 25:18]
  reg [31:0] _RAND_20;
  reg [15:0] gamma_1_7; // @[Frontend.scala 25:18]
  reg [31:0] _RAND_21;
  reg [15:0] gamma_2_0; // @[Frontend.scala 25:18]
  reg [31:0] _RAND_22;
  reg [15:0] gamma_2_1; // @[Frontend.scala 25:18]
  reg [31:0] _RAND_23;
  reg [15:0] gamma_2_2; // @[Frontend.scala 25:18]
  reg [31:0] _RAND_24;
  reg [15:0] gamma_2_3; // @[Frontend.scala 25:18]
  reg [31:0] _RAND_25;
  reg [15:0] gamma_2_4; // @[Frontend.scala 25:18]
  reg [31:0] _RAND_26;
  reg [15:0] gamma_2_5; // @[Frontend.scala 25:18]
  reg [31:0] _RAND_27;
  reg [15:0] gamma_2_6; // @[Frontend.scala 25:18]
  reg [31:0] _RAND_28;
  reg [15:0] gamma_2_7; // @[Frontend.scala 25:18]
  reg [31:0] _RAND_29;
  reg [15:0] gamma_3_0; // @[Frontend.scala 25:18]
  reg [31:0] _RAND_30;
  reg [15:0] gamma_3_1; // @[Frontend.scala 25:18]
  reg [31:0] _RAND_31;
  reg [15:0] gamma_3_2; // @[Frontend.scala 25:18]
  reg [31:0] _RAND_32;
  reg [15:0] gamma_3_3; // @[Frontend.scala 25:18]
  reg [31:0] _RAND_33;
  reg [15:0] gamma_3_4; // @[Frontend.scala 25:18]
  reg [31:0] _RAND_34;
  reg [15:0] gamma_3_5; // @[Frontend.scala 25:18]
  reg [31:0] _RAND_35;
  reg [15:0] gamma_3_6; // @[Frontend.scala 25:18]
  reg [31:0] _RAND_36;
  reg [15:0] gamma_3_7; // @[Frontend.scala 25:18]
  reg [31:0] _RAND_37;
  reg [15:0] localWeights_0_0; // @[Frontend.scala 27:25]
  reg [31:0] _RAND_38;
  reg [15:0] localWeights_0_1; // @[Frontend.scala 27:25]
  reg [31:0] _RAND_39;
  reg [15:0] localWeights_0_2; // @[Frontend.scala 27:25]
  reg [31:0] _RAND_40;
  reg [15:0] localWeights_0_3; // @[Frontend.scala 27:25]
  reg [31:0] _RAND_41;
  reg [15:0] localWeights_0_4; // @[Frontend.scala 27:25]
  reg [31:0] _RAND_42;
  reg [15:0] localWeights_0_5; // @[Frontend.scala 27:25]
  reg [31:0] _RAND_43;
  reg [15:0] localWeights_0_6; // @[Frontend.scala 27:25]
  reg [31:0] _RAND_44;
  reg [15:0] localWeights_0_7; // @[Frontend.scala 27:25]
  reg [31:0] _RAND_45;
  reg [15:0] localWeights_1_0; // @[Frontend.scala 27:25]
  reg [31:0] _RAND_46;
  reg [15:0] localWeights_1_1; // @[Frontend.scala 27:25]
  reg [31:0] _RAND_47;
  reg [15:0] localWeights_1_2; // @[Frontend.scala 27:25]
  reg [31:0] _RAND_48;
  reg [15:0] localWeights_1_3; // @[Frontend.scala 27:25]
  reg [31:0] _RAND_49;
  reg [15:0] localWeights_1_4; // @[Frontend.scala 27:25]
  reg [31:0] _RAND_50;
  reg [15:0] localWeights_1_5; // @[Frontend.scala 27:25]
  reg [31:0] _RAND_51;
  reg [15:0] localWeights_1_6; // @[Frontend.scala 27:25]
  reg [31:0] _RAND_52;
  reg [15:0] localWeights_1_7; // @[Frontend.scala 27:25]
  reg [31:0] _RAND_53;
  reg [15:0] localWeights_2_0; // @[Frontend.scala 27:25]
  reg [31:0] _RAND_54;
  reg [15:0] localWeights_2_1; // @[Frontend.scala 27:25]
  reg [31:0] _RAND_55;
  reg [15:0] localWeights_2_2; // @[Frontend.scala 27:25]
  reg [31:0] _RAND_56;
  reg [15:0] localWeights_2_3; // @[Frontend.scala 27:25]
  reg [31:0] _RAND_57;
  reg [15:0] localWeights_2_4; // @[Frontend.scala 27:25]
  reg [31:0] _RAND_58;
  reg [15:0] localWeights_2_5; // @[Frontend.scala 27:25]
  reg [31:0] _RAND_59;
  reg [15:0] localWeights_2_6; // @[Frontend.scala 27:25]
  reg [31:0] _RAND_60;
  reg [15:0] localWeights_2_7; // @[Frontend.scala 27:25]
  reg [31:0] _RAND_61;
  reg [15:0] localWeights_3_0; // @[Frontend.scala 27:25]
  reg [31:0] _RAND_62;
  reg [15:0] localWeights_3_1; // @[Frontend.scala 27:25]
  reg [31:0] _RAND_63;
  reg [15:0] localWeights_3_2; // @[Frontend.scala 27:25]
  reg [31:0] _RAND_64;
  reg [15:0] localWeights_3_3; // @[Frontend.scala 27:25]
  reg [31:0] _RAND_65;
  reg [15:0] localWeights_3_4; // @[Frontend.scala 27:25]
  reg [31:0] _RAND_66;
  reg [15:0] localWeights_3_5; // @[Frontend.scala 27:25]
  reg [31:0] _RAND_67;
  reg [15:0] localWeights_3_6; // @[Frontend.scala 27:25]
  reg [31:0] _RAND_68;
  reg [15:0] localWeights_3_7; // @[Frontend.scala 27:25]
  reg [31:0] _RAND_69;
  wire  _T_6; // @[Frontend.scala 38:17]
  wire  _T_7; // @[Frontend.scala 42:19]
  wire [1:0] _T_9; // @[Frontend.scala 43:20]
  wire  _T_11; // @[Frontend.scala 52:27]
  wire  _T_12; // @[Frontend.scala 54:31]
  wire  _T_13; // @[Frontend.scala 54:28]
  wire  _T_14; // @[Frontend.scala 53:27]
  wire  _T_16; // @[Frontend.scala 55:28]
  wire  _T_17; // @[Frontend.scala 54:45]
  wire  _T_19; // @[Frontend.scala 56:29]
  wire  _T_20; // @[Frontend.scala 56:54]
  wire  _T_21; // @[Frontend.scala 56:45]
  wire  _T_22; // @[Frontend.scala 55:45]
  wire [15:0] _T_25; // @[Frontend.scala 63:42]
  wire [15:0] _T_27; // @[Frontend.scala 63:49]
  wire [15:0] _T_28; // @[Frontend.scala 63:49]
  wire [15:0] _T_29; // @[Frontend.scala 63:42]
  wire [15:0] _T_31; // @[Frontend.scala 63:49]
  wire [15:0] _T_32; // @[Frontend.scala 63:49]
  wire [15:0] _T_33; // @[Frontend.scala 63:42]
  wire [15:0] _T_35; // @[Frontend.scala 63:49]
  wire [15:0] _T_36; // @[Frontend.scala 63:49]
  wire [15:0] _T_37; // @[Frontend.scala 63:42]
  wire [15:0] _T_39; // @[Frontend.scala 63:49]
  wire [15:0] _T_40; // @[Frontend.scala 63:49]
  wire [15:0] _T_41; // @[Frontend.scala 63:42]
  wire [15:0] _T_43; // @[Frontend.scala 63:49]
  wire [15:0] _T_44; // @[Frontend.scala 63:49]
  wire [15:0] _T_45; // @[Frontend.scala 63:42]
  wire [15:0] _T_47; // @[Frontend.scala 63:49]
  wire [15:0] _T_48; // @[Frontend.scala 63:49]
  wire [15:0] _T_49; // @[Frontend.scala 63:42]
  wire [15:0] _T_51; // @[Frontend.scala 63:49]
  wire [15:0] _T_52; // @[Frontend.scala 63:49]
  wire [15:0] _T_53; // @[Frontend.scala 63:42]
  wire [15:0] _T_55; // @[Frontend.scala 63:49]
  wire [15:0] _T_56; // @[Frontend.scala 63:49]
  wire  _T_57; // @[Frontend.scala 65:23]
  wire [15:0] _T_58; // @[Frontend.scala 68:59]
  wire [15:0] _T_60; // @[Frontend.scala 68:42]
  wire [15:0] _T_61; // @[Frontend.scala 68:42]
  wire [15:0] _T_62; // @[Frontend.scala 68:59]
  wire [15:0] _T_64; // @[Frontend.scala 68:42]
  wire [15:0] _T_65; // @[Frontend.scala 68:42]
  wire [15:0] _T_66; // @[Frontend.scala 68:59]
  wire [15:0] _T_68; // @[Frontend.scala 68:42]
  wire [15:0] _T_69; // @[Frontend.scala 68:42]
  wire [15:0] _T_70; // @[Frontend.scala 68:59]
  wire [15:0] _T_72; // @[Frontend.scala 68:42]
  wire [15:0] _T_73; // @[Frontend.scala 68:42]
  wire [15:0] _T_74; // @[Frontend.scala 68:59]
  wire [15:0] _T_76; // @[Frontend.scala 68:42]
  wire [15:0] _T_77; // @[Frontend.scala 68:42]
  wire [15:0] _T_78; // @[Frontend.scala 68:59]
  wire [15:0] _T_80; // @[Frontend.scala 68:42]
  wire [15:0] _T_81; // @[Frontend.scala 68:42]
  wire [15:0] _T_82; // @[Frontend.scala 68:59]
  wire [15:0] _T_84; // @[Frontend.scala 68:42]
  wire [15:0] _T_85; // @[Frontend.scala 68:42]
  wire [15:0] _T_86; // @[Frontend.scala 68:59]
  wire [15:0] _T_88; // @[Frontend.scala 68:42]
  wire [15:0] _T_89; // @[Frontend.scala 68:42]
  wire [15:0] _GEN_70; // @[Frontend.scala 65:32]
  wire [15:0] _GEN_71; // @[Frontend.scala 65:32]
  wire [15:0] _GEN_72; // @[Frontend.scala 65:32]
  wire [15:0] _GEN_73; // @[Frontend.scala 65:32]
  wire [15:0] _GEN_74; // @[Frontend.scala 65:32]
  wire [15:0] _GEN_75; // @[Frontend.scala 65:32]
  wire [15:0] _GEN_76; // @[Frontend.scala 65:32]
  wire [15:0] _GEN_77; // @[Frontend.scala 65:32]
  wire [15:0] _GEN_118; // @[Frontend.scala 75:20]
  wire [15:0] _GEN_126; // @[Frontend.scala 75:20]
  wire [15:0] _GEN_134; // @[Frontend.scala 75:20]
  wire [15:0] _GEN_144; // @[Frontend.scala 58:28]
  wire [15:0] _GEN_119; // @[Frontend.scala 75:20]
  wire [15:0] _GEN_127; // @[Frontend.scala 75:20]
  wire [15:0] _GEN_135; // @[Frontend.scala 75:20]
  wire [15:0] _GEN_145; // @[Frontend.scala 58:28]
  wire [15:0] _GEN_120; // @[Frontend.scala 75:20]
  wire [15:0] _GEN_128; // @[Frontend.scala 75:20]
  wire [15:0] _GEN_136; // @[Frontend.scala 75:20]
  wire [15:0] _GEN_146; // @[Frontend.scala 58:28]
  wire [15:0] _GEN_121; // @[Frontend.scala 75:20]
  wire [15:0] _GEN_129; // @[Frontend.scala 75:20]
  wire [15:0] _GEN_137; // @[Frontend.scala 75:20]
  wire [15:0] _GEN_147; // @[Frontend.scala 58:28]
  wire [15:0] _GEN_122; // @[Frontend.scala 75:20]
  wire [15:0] _GEN_130; // @[Frontend.scala 75:20]
  wire [15:0] _GEN_138; // @[Frontend.scala 75:20]
  wire [15:0] _GEN_148; // @[Frontend.scala 58:28]
  wire [15:0] _GEN_123; // @[Frontend.scala 75:20]
  wire [15:0] _GEN_131; // @[Frontend.scala 75:20]
  wire [15:0] _GEN_139; // @[Frontend.scala 75:20]
  wire [15:0] _GEN_149; // @[Frontend.scala 58:28]
  wire [15:0] _GEN_124; // @[Frontend.scala 75:20]
  wire [15:0] _GEN_132; // @[Frontend.scala 75:20]
  wire [15:0] _GEN_140; // @[Frontend.scala 75:20]
  wire [15:0] _GEN_150; // @[Frontend.scala 58:28]
  wire [15:0] _GEN_125; // @[Frontend.scala 75:20]
  wire [15:0] _GEN_133; // @[Frontend.scala 75:20]
  wire [15:0] _GEN_141; // @[Frontend.scala 75:20]
  wire [15:0] _GEN_151; // @[Frontend.scala 58:28]
  wire  _GEN_143; // @[Frontend.scala 58:28]
  wire [1:0] _T_90; // @[Frontend.scala 80:23]
  wire [4:0] _T_91; // @[Frontend.scala 81:23]
  wire [2:0] _T_92;
  wire  _GEN_497; // @[Frontend.scala 82:31]
  wire  _GEN_498; // @[Frontend.scala 82:31]
  wire [15:0] _GEN_185; // @[Frontend.scala 82:31]
  wire  _GEN_500; // @[Frontend.scala 82:31]
  wire [15:0] _GEN_186; // @[Frontend.scala 82:31]
  wire  _GEN_502; // @[Frontend.scala 82:31]
  wire [15:0] _GEN_187; // @[Frontend.scala 82:31]
  wire  _GEN_504; // @[Frontend.scala 82:31]
  wire [15:0] _GEN_188; // @[Frontend.scala 82:31]
  wire  _GEN_506; // @[Frontend.scala 82:31]
  wire [15:0] _GEN_189; // @[Frontend.scala 82:31]
  wire  _GEN_508; // @[Frontend.scala 82:31]
  wire [15:0] _GEN_190; // @[Frontend.scala 82:31]
  wire  _GEN_510; // @[Frontend.scala 82:31]
  wire [15:0] _GEN_191; // @[Frontend.scala 82:31]
  wire  _GEN_511; // @[Frontend.scala 82:31]
  wire  _GEN_512; // @[Frontend.scala 82:31]
  wire [15:0] _GEN_192; // @[Frontend.scala 82:31]
  wire [15:0] _GEN_193; // @[Frontend.scala 82:31]
  wire [15:0] _GEN_194; // @[Frontend.scala 82:31]
  wire [15:0] _GEN_195; // @[Frontend.scala 82:31]
  wire [15:0] _GEN_196; // @[Frontend.scala 82:31]
  wire [15:0] _GEN_197; // @[Frontend.scala 82:31]
  wire [15:0] _GEN_198; // @[Frontend.scala 82:31]
  wire [15:0] _GEN_199; // @[Frontend.scala 82:31]
  wire  _GEN_527; // @[Frontend.scala 82:31]
  wire [15:0] _GEN_200; // @[Frontend.scala 82:31]
  wire [15:0] _GEN_201; // @[Frontend.scala 82:31]
  wire [15:0] _GEN_202; // @[Frontend.scala 82:31]
  wire [15:0] _GEN_203; // @[Frontend.scala 82:31]
  wire [15:0] _GEN_204; // @[Frontend.scala 82:31]
  wire [15:0] _GEN_205; // @[Frontend.scala 82:31]
  wire [15:0] _GEN_206; // @[Frontend.scala 82:31]
  wire [15:0] _GEN_207; // @[Frontend.scala 82:31]
  wire  _GEN_543; // @[Frontend.scala 82:31]
  wire [15:0] _GEN_208; // @[Frontend.scala 82:31]
  wire [15:0] _GEN_209; // @[Frontend.scala 82:31]
  wire [15:0] _GEN_210; // @[Frontend.scala 82:31]
  wire [15:0] _GEN_211; // @[Frontend.scala 82:31]
  wire [15:0] _GEN_212; // @[Frontend.scala 82:31]
  wire [15:0] _GEN_213; // @[Frontend.scala 82:31]
  wire [15:0] _GEN_214; // @[Frontend.scala 82:31]
  wire [15:0] _GEN_215; // @[Frontend.scala 82:31]
  wire [15:0] _T_93; // @[Frontend.scala 82:31]
  wire [31:0] _T_94; // @[Frontend.scala 84:33]
  wire [21:0] _T_95; // @[Frontend.scala 84:47]
  wire [15:0] _T_96; // @[Frontend.scala 84:78]
  wire [21:0] _GEN_559; // @[Frontend.scala 84:61]
  wire [21:0] _T_98; // @[Frontend.scala 84:61]
  wire [21:0] _T_99; // @[Frontend.scala 84:61]
  wire [31:0] _T_100; // @[Frontend.scala 84:33]
  wire [21:0] _T_101; // @[Frontend.scala 84:47]
  wire [15:0] _T_102; // @[Frontend.scala 84:78]
  wire [21:0] _GEN_560; // @[Frontend.scala 84:61]
  wire [21:0] _T_104; // @[Frontend.scala 84:61]
  wire [21:0] _T_105; // @[Frontend.scala 84:61]
  wire [31:0] _T_106; // @[Frontend.scala 84:33]
  wire [21:0] _T_107; // @[Frontend.scala 84:47]
  wire [15:0] _T_108; // @[Frontend.scala 84:78]
  wire [21:0] _GEN_561; // @[Frontend.scala 84:61]
  wire [21:0] _T_110; // @[Frontend.scala 84:61]
  wire [21:0] _T_111; // @[Frontend.scala 84:61]
  wire [31:0] _T_112; // @[Frontend.scala 84:33]
  wire [21:0] _T_113; // @[Frontend.scala 84:47]
  wire [15:0] _T_114; // @[Frontend.scala 84:78]
  wire [21:0] _GEN_562; // @[Frontend.scala 84:61]
  wire [21:0] _T_116; // @[Frontend.scala 84:61]
  wire [21:0] _T_117; // @[Frontend.scala 84:61]
  wire [31:0] _T_118; // @[Frontend.scala 84:33]
  wire [21:0] _T_119; // @[Frontend.scala 84:47]
  wire [15:0] _T_120; // @[Frontend.scala 84:78]
  wire [21:0] _GEN_563; // @[Frontend.scala 84:61]
  wire [21:0] _T_122; // @[Frontend.scala 84:61]
  wire [21:0] _T_123; // @[Frontend.scala 84:61]
  wire [31:0] _T_124; // @[Frontend.scala 84:33]
  wire [21:0] _T_125; // @[Frontend.scala 84:47]
  wire [15:0] _T_126; // @[Frontend.scala 84:78]
  wire [21:0] _GEN_564; // @[Frontend.scala 84:61]
  wire [21:0] _T_128; // @[Frontend.scala 84:61]
  wire [21:0] _T_129; // @[Frontend.scala 84:61]
  wire [31:0] _T_130; // @[Frontend.scala 84:33]
  wire [21:0] _T_131; // @[Frontend.scala 84:47]
  wire [15:0] _T_132; // @[Frontend.scala 84:78]
  wire [21:0] _GEN_565; // @[Frontend.scala 84:61]
  wire [21:0] _T_134; // @[Frontend.scala 84:61]
  wire [21:0] _T_135; // @[Frontend.scala 84:61]
  wire [31:0] _T_136; // @[Frontend.scala 84:33]
  wire [21:0] _T_137; // @[Frontend.scala 84:47]
  wire [15:0] _T_138; // @[Frontend.scala 84:78]
  wire [21:0] _GEN_566; // @[Frontend.scala 84:61]
  wire [21:0] _T_140; // @[Frontend.scala 84:61]
  wire [21:0] _T_141; // @[Frontend.scala 84:61]
  wire  _T_142; // @[SliceCounter.scala 22:15]
  wire [1:0] _T_144; // @[SliceCounter.scala 23:16]
  wire  _T_145; // @[SliceCounter.scala 26:16]
  wire [4:0] _T_147; // @[SliceCounter.scala 27:16]
  wire  _T_148; // @[SliceCounter.scala 31:18]
  wire [4:0] _T_150; // @[SliceCounter.scala 32:18]
  wire [4:0] _T_152; // @[SliceCounter.scala 33:18]
  wire  _GEN_231; // @[Frontend.scala 56:64]
  wire  _GEN_232; // @[Frontend.scala 56:64]
  wire  _GEN_280; // @[Frontend.scala 49:34]
  wire  _GEN_281; // @[Frontend.scala 49:34]
  wire  _GEN_314; // @[Frontend.scala 49:34]
  wire  _GEN_329; // @[Frontend.scala 38:26]
  wire  _GEN_364; // @[Frontend.scala 38:26]
  wire  _GEN_365; // @[Frontend.scala 38:26]
  wire  _GEN_398; // @[Frontend.scala 38:26]
  wire [15:0] _GEN_567; // @[Frontend.scala 84:26]
  wire [15:0] _GEN_568; // @[Frontend.scala 84:26]
  wire [15:0] _GEN_569; // @[Frontend.scala 84:26]
  wire [15:0] _GEN_570; // @[Frontend.scala 84:26]
  wire [15:0] _GEN_571; // @[Frontend.scala 84:26]
  wire [15:0] _GEN_572; // @[Frontend.scala 84:26]
  wire [15:0] _GEN_573; // @[Frontend.scala 84:26]
  wire [15:0] _GEN_574; // @[Frontend.scala 84:26]
  assign _T_6 = phase == 1'h0; // @[Frontend.scala 38:17]
  assign _T_7 = jj != 2'h2; // @[Frontend.scala 42:19]
  assign _T_9 = jj + 2'h1; // @[Frontend.scala 43:20]
  assign _T_11 = io_off_ready & io_mi1_valid; // @[Frontend.scala 52:27]
  assign _T_12 = _T_5 == 1'h0; // @[Frontend.scala 54:31]
  assign _T_13 = io_a0_valid | _T_12; // @[Frontend.scala 54:28]
  assign _T_14 = _T_11 & _T_13; // @[Frontend.scala 53:27]
  assign _T_16 = io_wi_valid | _T_12; // @[Frontend.scala 55:28]
  assign _T_17 = _T_14 & _T_16; // @[Frontend.scala 54:45]
  assign _T_19 = io_adj_valid | _T_12; // @[Frontend.scala 56:29]
  assign _T_20 = _T_2 == 5'h0; // @[Frontend.scala 56:54]
  assign _T_21 = _T_19 | _T_20; // @[Frontend.scala 56:45]
  assign _T_22 = _T_17 & _T_21; // @[Frontend.scala 55:45]
  assign _T_25 = $signed(io_a0_bits_0); // @[Frontend.scala 63:42]
  assign _T_27 = $signed(_T_25) + $signed(io_wi_bits_0); // @[Frontend.scala 63:49]
  assign _T_28 = $signed(_T_27); // @[Frontend.scala 63:49]
  assign _T_29 = $signed(io_a0_bits_1); // @[Frontend.scala 63:42]
  assign _T_31 = $signed(_T_29) + $signed(io_wi_bits_1); // @[Frontend.scala 63:49]
  assign _T_32 = $signed(_T_31); // @[Frontend.scala 63:49]
  assign _T_33 = $signed(io_a0_bits_2); // @[Frontend.scala 63:42]
  assign _T_35 = $signed(_T_33) + $signed(io_wi_bits_2); // @[Frontend.scala 63:49]
  assign _T_36 = $signed(_T_35); // @[Frontend.scala 63:49]
  assign _T_37 = $signed(io_a0_bits_3); // @[Frontend.scala 63:42]
  assign _T_39 = $signed(_T_37) + $signed(io_wi_bits_3); // @[Frontend.scala 63:49]
  assign _T_40 = $signed(_T_39); // @[Frontend.scala 63:49]
  assign _T_41 = $signed(io_a0_bits_4); // @[Frontend.scala 63:42]
  assign _T_43 = $signed(_T_41) + $signed(io_wi_bits_4); // @[Frontend.scala 63:49]
  assign _T_44 = $signed(_T_43); // @[Frontend.scala 63:49]
  assign _T_45 = $signed(io_a0_bits_5); // @[Frontend.scala 63:42]
  assign _T_47 = $signed(_T_45) + $signed(io_wi_bits_5); // @[Frontend.scala 63:49]
  assign _T_48 = $signed(_T_47); // @[Frontend.scala 63:49]
  assign _T_49 = $signed(io_a0_bits_6); // @[Frontend.scala 63:42]
  assign _T_51 = $signed(_T_49) + $signed(io_wi_bits_6); // @[Frontend.scala 63:49]
  assign _T_52 = $signed(_T_51); // @[Frontend.scala 63:49]
  assign _T_53 = $signed(io_a0_bits_7); // @[Frontend.scala 63:42]
  assign _T_55 = $signed(_T_53) + $signed(io_wi_bits_7); // @[Frontend.scala 63:49]
  assign _T_56 = $signed(_T_55); // @[Frontend.scala 63:49]
  assign _T_57 = _T_2 != 5'h0; // @[Frontend.scala 65:23]
  assign _T_58 = $signed(io_adj_bits_0); // @[Frontend.scala 68:59]
  assign _T_60 = $signed(_T_28) + $signed(_T_58); // @[Frontend.scala 68:42]
  assign _T_61 = $signed(_T_60); // @[Frontend.scala 68:42]
  assign _T_62 = $signed(io_adj_bits_1); // @[Frontend.scala 68:59]
  assign _T_64 = $signed(_T_32) + $signed(_T_62); // @[Frontend.scala 68:42]
  assign _T_65 = $signed(_T_64); // @[Frontend.scala 68:42]
  assign _T_66 = $signed(io_adj_bits_2); // @[Frontend.scala 68:59]
  assign _T_68 = $signed(_T_36) + $signed(_T_66); // @[Frontend.scala 68:42]
  assign _T_69 = $signed(_T_68); // @[Frontend.scala 68:42]
  assign _T_70 = $signed(io_adj_bits_3); // @[Frontend.scala 68:59]
  assign _T_72 = $signed(_T_40) + $signed(_T_70); // @[Frontend.scala 68:42]
  assign _T_73 = $signed(_T_72); // @[Frontend.scala 68:42]
  assign _T_74 = $signed(io_adj_bits_4); // @[Frontend.scala 68:59]
  assign _T_76 = $signed(_T_44) + $signed(_T_74); // @[Frontend.scala 68:42]
  assign _T_77 = $signed(_T_76); // @[Frontend.scala 68:42]
  assign _T_78 = $signed(io_adj_bits_5); // @[Frontend.scala 68:59]
  assign _T_80 = $signed(_T_48) + $signed(_T_78); // @[Frontend.scala 68:42]
  assign _T_81 = $signed(_T_80); // @[Frontend.scala 68:42]
  assign _T_82 = $signed(io_adj_bits_6); // @[Frontend.scala 68:59]
  assign _T_84 = $signed(_T_52) + $signed(_T_82); // @[Frontend.scala 68:42]
  assign _T_85 = $signed(_T_84); // @[Frontend.scala 68:42]
  assign _T_86 = $signed(io_adj_bits_7); // @[Frontend.scala 68:59]
  assign _T_88 = $signed(_T_56) + $signed(_T_86); // @[Frontend.scala 68:42]
  assign _T_89 = $signed(_T_88); // @[Frontend.scala 68:42]
  assign _GEN_70 = _T_57 ? $signed(_T_61) : $signed(_T_28); // @[Frontend.scala 65:32]
  assign _GEN_71 = _T_57 ? $signed(_T_65) : $signed(_T_32); // @[Frontend.scala 65:32]
  assign _GEN_72 = _T_57 ? $signed(_T_69) : $signed(_T_36); // @[Frontend.scala 65:32]
  assign _GEN_73 = _T_57 ? $signed(_T_73) : $signed(_T_40); // @[Frontend.scala 65:32]
  assign _GEN_74 = _T_57 ? $signed(_T_77) : $signed(_T_44); // @[Frontend.scala 65:32]
  assign _GEN_75 = _T_57 ? $signed(_T_81) : $signed(_T_48); // @[Frontend.scala 65:32]
  assign _GEN_76 = _T_57 ? $signed(_T_85) : $signed(_T_52); // @[Frontend.scala 65:32]
  assign _GEN_77 = _T_57 ? $signed(_T_89) : $signed(_T_56); // @[Frontend.scala 65:32]
  assign _GEN_118 = 2'h1 == _T ? $signed(localWeights_1_0) : $signed(localWeights_0_0); // @[Frontend.scala 75:20]
  assign _GEN_126 = 2'h2 == _T ? $signed(localWeights_2_0) : $signed(_GEN_118); // @[Frontend.scala 75:20]
  assign _GEN_134 = 2'h3 == _T ? $signed(localWeights_3_0) : $signed(_GEN_126); // @[Frontend.scala 75:20]
  assign _GEN_144 = _T_5 ? $signed(_GEN_70) : $signed(_GEN_134); // @[Frontend.scala 58:28]
  assign _GEN_119 = 2'h1 == _T ? $signed(localWeights_1_1) : $signed(localWeights_0_1); // @[Frontend.scala 75:20]
  assign _GEN_127 = 2'h2 == _T ? $signed(localWeights_2_1) : $signed(_GEN_119); // @[Frontend.scala 75:20]
  assign _GEN_135 = 2'h3 == _T ? $signed(localWeights_3_1) : $signed(_GEN_127); // @[Frontend.scala 75:20]
  assign _GEN_145 = _T_5 ? $signed(_GEN_71) : $signed(_GEN_135); // @[Frontend.scala 58:28]
  assign _GEN_120 = 2'h1 == _T ? $signed(localWeights_1_2) : $signed(localWeights_0_2); // @[Frontend.scala 75:20]
  assign _GEN_128 = 2'h2 == _T ? $signed(localWeights_2_2) : $signed(_GEN_120); // @[Frontend.scala 75:20]
  assign _GEN_136 = 2'h3 == _T ? $signed(localWeights_3_2) : $signed(_GEN_128); // @[Frontend.scala 75:20]
  assign _GEN_146 = _T_5 ? $signed(_GEN_72) : $signed(_GEN_136); // @[Frontend.scala 58:28]
  assign _GEN_121 = 2'h1 == _T ? $signed(localWeights_1_3) : $signed(localWeights_0_3); // @[Frontend.scala 75:20]
  assign _GEN_129 = 2'h2 == _T ? $signed(localWeights_2_3) : $signed(_GEN_121); // @[Frontend.scala 75:20]
  assign _GEN_137 = 2'h3 == _T ? $signed(localWeights_3_3) : $signed(_GEN_129); // @[Frontend.scala 75:20]
  assign _GEN_147 = _T_5 ? $signed(_GEN_73) : $signed(_GEN_137); // @[Frontend.scala 58:28]
  assign _GEN_122 = 2'h1 == _T ? $signed(localWeights_1_4) : $signed(localWeights_0_4); // @[Frontend.scala 75:20]
  assign _GEN_130 = 2'h2 == _T ? $signed(localWeights_2_4) : $signed(_GEN_122); // @[Frontend.scala 75:20]
  assign _GEN_138 = 2'h3 == _T ? $signed(localWeights_3_4) : $signed(_GEN_130); // @[Frontend.scala 75:20]
  assign _GEN_148 = _T_5 ? $signed(_GEN_74) : $signed(_GEN_138); // @[Frontend.scala 58:28]
  assign _GEN_123 = 2'h1 == _T ? $signed(localWeights_1_5) : $signed(localWeights_0_5); // @[Frontend.scala 75:20]
  assign _GEN_131 = 2'h2 == _T ? $signed(localWeights_2_5) : $signed(_GEN_123); // @[Frontend.scala 75:20]
  assign _GEN_139 = 2'h3 == _T ? $signed(localWeights_3_5) : $signed(_GEN_131); // @[Frontend.scala 75:20]
  assign _GEN_149 = _T_5 ? $signed(_GEN_75) : $signed(_GEN_139); // @[Frontend.scala 58:28]
  assign _GEN_124 = 2'h1 == _T ? $signed(localWeights_1_6) : $signed(localWeights_0_6); // @[Frontend.scala 75:20]
  assign _GEN_132 = 2'h2 == _T ? $signed(localWeights_2_6) : $signed(_GEN_124); // @[Frontend.scala 75:20]
  assign _GEN_140 = 2'h3 == _T ? $signed(localWeights_3_6) : $signed(_GEN_132); // @[Frontend.scala 75:20]
  assign _GEN_150 = _T_5 ? $signed(_GEN_76) : $signed(_GEN_140); // @[Frontend.scala 58:28]
  assign _GEN_125 = 2'h1 == _T ? $signed(localWeights_1_7) : $signed(localWeights_0_7); // @[Frontend.scala 75:20]
  assign _GEN_133 = 2'h2 == _T ? $signed(localWeights_2_7) : $signed(_GEN_125); // @[Frontend.scala 75:20]
  assign _GEN_141 = 2'h3 == _T ? $signed(localWeights_3_7) : $signed(_GEN_133); // @[Frontend.scala 75:20]
  assign _GEN_151 = _T_5 ? $signed(_GEN_77) : $signed(_GEN_141); // @[Frontend.scala 58:28]
  assign _GEN_143 = _T_5 ? _T_57 : 1'h0; // @[Frontend.scala 58:28]
  assign _T_90 = _T_1[4:3]; // @[Frontend.scala 80:23]
  assign _T_91 = _T_1 & 5'h7; // @[Frontend.scala 81:23]
  assign _T_92 = _T_91[2:0];
  assign _GEN_497 = 2'h0 == _T_90; // @[Frontend.scala 82:31]
  assign _GEN_498 = 3'h1 == _T_92; // @[Frontend.scala 82:31]
  assign _GEN_185 = _GEN_497 & _GEN_498 ? gamma_0_1 : gamma_0_0; // @[Frontend.scala 82:31]
  assign _GEN_500 = 3'h2 == _T_92; // @[Frontend.scala 82:31]
  assign _GEN_186 = _GEN_497 & _GEN_500 ? gamma_0_2 : _GEN_185; // @[Frontend.scala 82:31]
  assign _GEN_502 = 3'h3 == _T_92; // @[Frontend.scala 82:31]
  assign _GEN_187 = _GEN_497 & _GEN_502 ? gamma_0_3 : _GEN_186; // @[Frontend.scala 82:31]
  assign _GEN_504 = 3'h4 == _T_92; // @[Frontend.scala 82:31]
  assign _GEN_188 = _GEN_497 & _GEN_504 ? gamma_0_4 : _GEN_187; // @[Frontend.scala 82:31]
  assign _GEN_506 = 3'h5 == _T_92; // @[Frontend.scala 82:31]
  assign _GEN_189 = _GEN_497 & _GEN_506 ? gamma_0_5 : _GEN_188; // @[Frontend.scala 82:31]
  assign _GEN_508 = 3'h6 == _T_92; // @[Frontend.scala 82:31]
  assign _GEN_190 = _GEN_497 & _GEN_508 ? gamma_0_6 : _GEN_189; // @[Frontend.scala 82:31]
  assign _GEN_510 = 3'h7 == _T_92; // @[Frontend.scala 82:31]
  assign _GEN_191 = _GEN_497 & _GEN_510 ? gamma_0_7 : _GEN_190; // @[Frontend.scala 82:31]
  assign _GEN_511 = 2'h1 == _T_90; // @[Frontend.scala 82:31]
  assign _GEN_512 = 3'h0 == _T_92; // @[Frontend.scala 82:31]
  assign _GEN_192 = _GEN_511 & _GEN_512 ? gamma_1_0 : _GEN_191; // @[Frontend.scala 82:31]
  assign _GEN_193 = _GEN_511 & _GEN_498 ? gamma_1_1 : _GEN_192; // @[Frontend.scala 82:31]
  assign _GEN_194 = _GEN_511 & _GEN_500 ? gamma_1_2 : _GEN_193; // @[Frontend.scala 82:31]
  assign _GEN_195 = _GEN_511 & _GEN_502 ? gamma_1_3 : _GEN_194; // @[Frontend.scala 82:31]
  assign _GEN_196 = _GEN_511 & _GEN_504 ? gamma_1_4 : _GEN_195; // @[Frontend.scala 82:31]
  assign _GEN_197 = _GEN_511 & _GEN_506 ? gamma_1_5 : _GEN_196; // @[Frontend.scala 82:31]
  assign _GEN_198 = _GEN_511 & _GEN_508 ? gamma_1_6 : _GEN_197; // @[Frontend.scala 82:31]
  assign _GEN_199 = _GEN_511 & _GEN_510 ? gamma_1_7 : _GEN_198; // @[Frontend.scala 82:31]
  assign _GEN_527 = 2'h2 == _T_90; // @[Frontend.scala 82:31]
  assign _GEN_200 = _GEN_527 & _GEN_512 ? gamma_2_0 : _GEN_199; // @[Frontend.scala 82:31]
  assign _GEN_201 = _GEN_527 & _GEN_498 ? gamma_2_1 : _GEN_200; // @[Frontend.scala 82:31]
  assign _GEN_202 = _GEN_527 & _GEN_500 ? gamma_2_2 : _GEN_201; // @[Frontend.scala 82:31]
  assign _GEN_203 = _GEN_527 & _GEN_502 ? gamma_2_3 : _GEN_202; // @[Frontend.scala 82:31]
  assign _GEN_204 = _GEN_527 & _GEN_504 ? gamma_2_4 : _GEN_203; // @[Frontend.scala 82:31]
  assign _GEN_205 = _GEN_527 & _GEN_506 ? gamma_2_5 : _GEN_204; // @[Frontend.scala 82:31]
  assign _GEN_206 = _GEN_527 & _GEN_508 ? gamma_2_6 : _GEN_205; // @[Frontend.scala 82:31]
  assign _GEN_207 = _GEN_527 & _GEN_510 ? gamma_2_7 : _GEN_206; // @[Frontend.scala 82:31]
  assign _GEN_543 = 2'h3 == _T_90; // @[Frontend.scala 82:31]
  assign _GEN_208 = _GEN_543 & _GEN_512 ? gamma_3_0 : _GEN_207; // @[Frontend.scala 82:31]
  assign _GEN_209 = _GEN_543 & _GEN_498 ? gamma_3_1 : _GEN_208; // @[Frontend.scala 82:31]
  assign _GEN_210 = _GEN_543 & _GEN_500 ? gamma_3_2 : _GEN_209; // @[Frontend.scala 82:31]
  assign _GEN_211 = _GEN_543 & _GEN_502 ? gamma_3_3 : _GEN_210; // @[Frontend.scala 82:31]
  assign _GEN_212 = _GEN_543 & _GEN_504 ? gamma_3_4 : _GEN_211; // @[Frontend.scala 82:31]
  assign _GEN_213 = _GEN_543 & _GEN_506 ? gamma_3_5 : _GEN_212; // @[Frontend.scala 82:31]
  assign _GEN_214 = _GEN_543 & _GEN_508 ? gamma_3_6 : _GEN_213; // @[Frontend.scala 82:31]
  assign _GEN_215 = _GEN_543 & _GEN_510 ? gamma_3_7 : _GEN_214; // @[Frontend.scala 82:31]
  assign _T_93 = $signed(_GEN_215); // @[Frontend.scala 82:31]
  assign _T_94 = $signed(_T_93) * $signed(_GEN_144); // @[Frontend.scala 84:33]
  assign _T_95 = _T_94[31:10]; // @[Frontend.scala 84:47]
  assign _T_96 = $signed(io_mi1_bits_0); // @[Frontend.scala 84:78]
  assign _GEN_559 = {{6{_T_96[15]}},_T_96}; // @[Frontend.scala 84:61]
  assign _T_98 = $signed(_T_95) - $signed(_GEN_559); // @[Frontend.scala 84:61]
  assign _T_99 = $signed(_T_98); // @[Frontend.scala 84:61]
  assign _T_100 = $signed(_T_93) * $signed(_GEN_145); // @[Frontend.scala 84:33]
  assign _T_101 = _T_100[31:10]; // @[Frontend.scala 84:47]
  assign _T_102 = $signed(io_mi1_bits_1); // @[Frontend.scala 84:78]
  assign _GEN_560 = {{6{_T_102[15]}},_T_102}; // @[Frontend.scala 84:61]
  assign _T_104 = $signed(_T_101) - $signed(_GEN_560); // @[Frontend.scala 84:61]
  assign _T_105 = $signed(_T_104); // @[Frontend.scala 84:61]
  assign _T_106 = $signed(_T_93) * $signed(_GEN_146); // @[Frontend.scala 84:33]
  assign _T_107 = _T_106[31:10]; // @[Frontend.scala 84:47]
  assign _T_108 = $signed(io_mi1_bits_2); // @[Frontend.scala 84:78]
  assign _GEN_561 = {{6{_T_108[15]}},_T_108}; // @[Frontend.scala 84:61]
  assign _T_110 = $signed(_T_107) - $signed(_GEN_561); // @[Frontend.scala 84:61]
  assign _T_111 = $signed(_T_110); // @[Frontend.scala 84:61]
  assign _T_112 = $signed(_T_93) * $signed(_GEN_147); // @[Frontend.scala 84:33]
  assign _T_113 = _T_112[31:10]; // @[Frontend.scala 84:47]
  assign _T_114 = $signed(io_mi1_bits_3); // @[Frontend.scala 84:78]
  assign _GEN_562 = {{6{_T_114[15]}},_T_114}; // @[Frontend.scala 84:61]
  assign _T_116 = $signed(_T_113) - $signed(_GEN_562); // @[Frontend.scala 84:61]
  assign _T_117 = $signed(_T_116); // @[Frontend.scala 84:61]
  assign _T_118 = $signed(_T_93) * $signed(_GEN_148); // @[Frontend.scala 84:33]
  assign _T_119 = _T_118[31:10]; // @[Frontend.scala 84:47]
  assign _T_120 = $signed(io_mi1_bits_4); // @[Frontend.scala 84:78]
  assign _GEN_563 = {{6{_T_120[15]}},_T_120}; // @[Frontend.scala 84:61]
  assign _T_122 = $signed(_T_119) - $signed(_GEN_563); // @[Frontend.scala 84:61]
  assign _T_123 = $signed(_T_122); // @[Frontend.scala 84:61]
  assign _T_124 = $signed(_T_93) * $signed(_GEN_149); // @[Frontend.scala 84:33]
  assign _T_125 = _T_124[31:10]; // @[Frontend.scala 84:47]
  assign _T_126 = $signed(io_mi1_bits_5); // @[Frontend.scala 84:78]
  assign _GEN_564 = {{6{_T_126[15]}},_T_126}; // @[Frontend.scala 84:61]
  assign _T_128 = $signed(_T_125) - $signed(_GEN_564); // @[Frontend.scala 84:61]
  assign _T_129 = $signed(_T_128); // @[Frontend.scala 84:61]
  assign _T_130 = $signed(_T_93) * $signed(_GEN_150); // @[Frontend.scala 84:33]
  assign _T_131 = _T_130[31:10]; // @[Frontend.scala 84:47]
  assign _T_132 = $signed(io_mi1_bits_6); // @[Frontend.scala 84:78]
  assign _GEN_565 = {{6{_T_132[15]}},_T_132}; // @[Frontend.scala 84:61]
  assign _T_134 = $signed(_T_131) - $signed(_GEN_565); // @[Frontend.scala 84:61]
  assign _T_135 = $signed(_T_134); // @[Frontend.scala 84:61]
  assign _T_136 = $signed(_T_93) * $signed(_GEN_151); // @[Frontend.scala 84:33]
  assign _T_137 = _T_136[31:10]; // @[Frontend.scala 84:47]
  assign _T_138 = $signed(io_mi1_bits_7); // @[Frontend.scala 84:78]
  assign _GEN_566 = {{6{_T_138[15]}},_T_138}; // @[Frontend.scala 84:61]
  assign _T_140 = $signed(_T_137) - $signed(_GEN_566); // @[Frontend.scala 84:61]
  assign _T_141 = $signed(_T_140); // @[Frontend.scala 84:61]
  assign _T_142 = _T != 2'h2; // @[SliceCounter.scala 22:15]
  assign _T_144 = _T + 2'h1; // @[SliceCounter.scala 23:16]
  assign _T_145 = _T_1 != 5'h17; // @[SliceCounter.scala 26:16]
  assign _T_147 = _T_1 + 5'h1; // @[SliceCounter.scala 27:16]
  assign _T_148 = _T_2 != 5'h16; // @[SliceCounter.scala 31:18]
  assign _T_150 = _T_2 + 5'h1; // @[SliceCounter.scala 32:18]
  assign _T_152 = _T_2 + 5'h2; // @[SliceCounter.scala 33:18]
  assign _GEN_231 = _T_22 ? _T_5 : 1'h0; // @[Frontend.scala 56:64]
  assign _GEN_232 = _T_22 ? _GEN_143 : 1'h0; // @[Frontend.scala 56:64]
  assign _GEN_280 = phase ? _GEN_231 : 1'h0; // @[Frontend.scala 49:34]
  assign _GEN_281 = phase ? _GEN_232 : 1'h0; // @[Frontend.scala 49:34]
  assign _GEN_314 = phase ? _T_22 : 1'h0; // @[Frontend.scala 49:34]
  assign _GEN_329 = _T_6 ? io_gi_valid : 1'h0; // @[Frontend.scala 38:26]
  assign _GEN_364 = _T_6 ? 1'h0 : _GEN_280; // @[Frontend.scala 38:26]
  assign _GEN_365 = _T_6 ? 1'h0 : _GEN_281; // @[Frontend.scala 38:26]
  assign _GEN_398 = _T_6 ? 1'h0 : _GEN_314; // @[Frontend.scala 38:26]
  assign io_gi_ready = io_start ? _GEN_329 : 1'h0; // @[Decoupled.scala 69:20 Frontend.scala 40:21]
  assign io_wi_ready = io_start ? _GEN_364 : 1'h0; // @[Decoupled.scala 69:20 Frontend.scala 61:23]
  assign io_a0_ready = io_start ? _GEN_364 : 1'h0; // @[Decoupled.scala 69:20 Frontend.scala 60:23]
  assign io_mi1_ready = io_start ? _GEN_398 : 1'h0; // @[Decoupled.scala 69:20 Frontend.scala 79:22]
  assign io_adj_ready = io_start ? _GEN_365 : 1'h0; // @[Decoupled.scala 69:20 Frontend.scala 66:26]
  assign io_off_valid = io_start ? _GEN_398 : 1'h0; // @[Decoupled.scala 53:20 Frontend.scala 78:22]
  assign _GEN_567 = _T_99[15:0]; // @[Frontend.scala 84:26]
  assign io_off_bits_0 = $signed(_GEN_567); // @[Frontend.scala 84:26]
  assign _GEN_568 = _T_105[15:0]; // @[Frontend.scala 84:26]
  assign io_off_bits_1 = $signed(_GEN_568); // @[Frontend.scala 84:26]
  assign _GEN_569 = _T_111[15:0]; // @[Frontend.scala 84:26]
  assign io_off_bits_2 = $signed(_GEN_569); // @[Frontend.scala 84:26]
  assign _GEN_570 = _T_117[15:0]; // @[Frontend.scala 84:26]
  assign io_off_bits_3 = $signed(_GEN_570); // @[Frontend.scala 84:26]
  assign _GEN_571 = _T_123[15:0]; // @[Frontend.scala 84:26]
  assign io_off_bits_4 = $signed(_GEN_571); // @[Frontend.scala 84:26]
  assign _GEN_572 = _T_129[15:0]; // @[Frontend.scala 84:26]
  assign io_off_bits_5 = $signed(_GEN_572); // @[Frontend.scala 84:26]
  assign _GEN_573 = _T_135[15:0]; // @[Frontend.scala 84:26]
  assign io_off_bits_6 = $signed(_GEN_573); // @[Frontend.scala 84:26]
  assign _GEN_574 = _T_141[15:0]; // @[Frontend.scala 84:26]
  assign io_off_bits_7 = $signed(_GEN_574); // @[Frontend.scala 84:26]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  phase = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  jj = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T = _RAND_2[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_1 = _RAND_3[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_2 = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_5 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  gamma_0_0 = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  gamma_0_1 = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  gamma_0_2 = _RAND_8[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  gamma_0_3 = _RAND_9[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  gamma_0_4 = _RAND_10[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  gamma_0_5 = _RAND_11[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  gamma_0_6 = _RAND_12[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  gamma_0_7 = _RAND_13[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  gamma_1_0 = _RAND_14[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  gamma_1_1 = _RAND_15[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  gamma_1_2 = _RAND_16[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  gamma_1_3 = _RAND_17[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  gamma_1_4 = _RAND_18[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  gamma_1_5 = _RAND_19[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  gamma_1_6 = _RAND_20[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  gamma_1_7 = _RAND_21[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  gamma_2_0 = _RAND_22[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  gamma_2_1 = _RAND_23[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  gamma_2_2 = _RAND_24[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  gamma_2_3 = _RAND_25[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  gamma_2_4 = _RAND_26[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  gamma_2_5 = _RAND_27[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  gamma_2_6 = _RAND_28[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  gamma_2_7 = _RAND_29[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  gamma_3_0 = _RAND_30[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  gamma_3_1 = _RAND_31[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  gamma_3_2 = _RAND_32[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  gamma_3_3 = _RAND_33[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  gamma_3_4 = _RAND_34[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  gamma_3_5 = _RAND_35[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  gamma_3_6 = _RAND_36[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  gamma_3_7 = _RAND_37[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  localWeights_0_0 = _RAND_38[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  localWeights_0_1 = _RAND_39[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  localWeights_0_2 = _RAND_40[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  localWeights_0_3 = _RAND_41[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  localWeights_0_4 = _RAND_42[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  localWeights_0_5 = _RAND_43[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  localWeights_0_6 = _RAND_44[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  localWeights_0_7 = _RAND_45[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  localWeights_1_0 = _RAND_46[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  localWeights_1_1 = _RAND_47[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  localWeights_1_2 = _RAND_48[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  localWeights_1_3 = _RAND_49[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  localWeights_1_4 = _RAND_50[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  localWeights_1_5 = _RAND_51[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  localWeights_1_6 = _RAND_52[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  localWeights_1_7 = _RAND_53[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  localWeights_2_0 = _RAND_54[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  localWeights_2_1 = _RAND_55[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  localWeights_2_2 = _RAND_56[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  localWeights_2_3 = _RAND_57[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  localWeights_2_4 = _RAND_58[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  localWeights_2_5 = _RAND_59[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  localWeights_2_6 = _RAND_60[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  localWeights_2_7 = _RAND_61[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  localWeights_3_0 = _RAND_62[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  localWeights_3_1 = _RAND_63[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  localWeights_3_2 = _RAND_64[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  localWeights_3_3 = _RAND_65[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  localWeights_3_4 = _RAND_66[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  localWeights_3_5 = _RAND_67[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  localWeights_3_6 = _RAND_68[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  localWeights_3_7 = _RAND_69[15:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      phase <= 1'h0;
    end else begin
      if (io_start) begin
        if (_T_6) begin
          if (io_gi_valid) begin
            if (!(_T_7)) begin
              phase <= 1'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      jj <= 2'h0;
    end else begin
      if (io_start) begin
        if (_T_6) begin
          if (io_gi_valid) begin
            if (_T_7) begin
              jj <= _T_9;
            end else begin
              jj <= 2'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      _T <= 2'h0;
    end else begin
      if (io_start) begin
        if (!(_T_6)) begin
          if (phase) begin
            if (_T_22) begin
              if (_T_142) begin
                _T <= _T_144;
              end else begin
                _T <= 2'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_1 <= 5'h1;
    end else begin
      if (io_start) begin
        if (!(_T_6)) begin
          if (phase) begin
            if (_T_22) begin
              if (!(_T_142)) begin
                if (_T_145) begin
                  _T_1 <= _T_147;
                end else begin
                  if (_T_148) begin
                    _T_1 <= _T_152;
                  end else begin
                    _T_1 <= 5'h1;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_2 <= 5'h0;
    end else begin
      if (io_start) begin
        if (!(_T_6)) begin
          if (phase) begin
            if (_T_22) begin
              if (!(_T_142)) begin
                if (!(_T_145)) begin
                  if (_T_148) begin
                    _T_2 <= _T_150;
                  end else begin
                    _T_2 <= 5'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_5 <= 1'h1;
    end else begin
      if (io_start) begin
        if (!(_T_6)) begin
          if (phase) begin
            if (_T_22) begin
              if (!(_T_142)) begin
                if (_T_145) begin
                  _T_5 <= 1'h0;
                end else begin
                  _T_5 <= 1'h1;
                end
              end
            end
          end
        end
      end
    end
    if (io_start) begin
      if (_T_6) begin
        if (io_gi_valid) begin
          if (2'h0 == jj) begin
            gamma_0_0 <= io_gi_bits_0;
          end
        end
      end
    end
    if (io_start) begin
      if (_T_6) begin
        if (io_gi_valid) begin
          if (2'h0 == jj) begin
            gamma_0_1 <= io_gi_bits_1;
          end
        end
      end
    end
    if (io_start) begin
      if (_T_6) begin
        if (io_gi_valid) begin
          if (2'h0 == jj) begin
            gamma_0_2 <= io_gi_bits_2;
          end
        end
      end
    end
    if (io_start) begin
      if (_T_6) begin
        if (io_gi_valid) begin
          if (2'h0 == jj) begin
            gamma_0_3 <= io_gi_bits_3;
          end
        end
      end
    end
    if (io_start) begin
      if (_T_6) begin
        if (io_gi_valid) begin
          if (2'h0 == jj) begin
            gamma_0_4 <= io_gi_bits_4;
          end
        end
      end
    end
    if (io_start) begin
      if (_T_6) begin
        if (io_gi_valid) begin
          if (2'h0 == jj) begin
            gamma_0_5 <= io_gi_bits_5;
          end
        end
      end
    end
    if (io_start) begin
      if (_T_6) begin
        if (io_gi_valid) begin
          if (2'h0 == jj) begin
            gamma_0_6 <= io_gi_bits_6;
          end
        end
      end
    end
    if (io_start) begin
      if (_T_6) begin
        if (io_gi_valid) begin
          if (2'h0 == jj) begin
            gamma_0_7 <= io_gi_bits_7;
          end
        end
      end
    end
    if (io_start) begin
      if (_T_6) begin
        if (io_gi_valid) begin
          if (2'h1 == jj) begin
            gamma_1_0 <= io_gi_bits_0;
          end
        end
      end
    end
    if (io_start) begin
      if (_T_6) begin
        if (io_gi_valid) begin
          if (2'h1 == jj) begin
            gamma_1_1 <= io_gi_bits_1;
          end
        end
      end
    end
    if (io_start) begin
      if (_T_6) begin
        if (io_gi_valid) begin
          if (2'h1 == jj) begin
            gamma_1_2 <= io_gi_bits_2;
          end
        end
      end
    end
    if (io_start) begin
      if (_T_6) begin
        if (io_gi_valid) begin
          if (2'h1 == jj) begin
            gamma_1_3 <= io_gi_bits_3;
          end
        end
      end
    end
    if (io_start) begin
      if (_T_6) begin
        if (io_gi_valid) begin
          if (2'h1 == jj) begin
            gamma_1_4 <= io_gi_bits_4;
          end
        end
      end
    end
    if (io_start) begin
      if (_T_6) begin
        if (io_gi_valid) begin
          if (2'h1 == jj) begin
            gamma_1_5 <= io_gi_bits_5;
          end
        end
      end
    end
    if (io_start) begin
      if (_T_6) begin
        if (io_gi_valid) begin
          if (2'h1 == jj) begin
            gamma_1_6 <= io_gi_bits_6;
          end
        end
      end
    end
    if (io_start) begin
      if (_T_6) begin
        if (io_gi_valid) begin
          if (2'h1 == jj) begin
            gamma_1_7 <= io_gi_bits_7;
          end
        end
      end
    end
    if (io_start) begin
      if (_T_6) begin
        if (io_gi_valid) begin
          if (2'h2 == jj) begin
            gamma_2_0 <= io_gi_bits_0;
          end
        end
      end
    end
    if (io_start) begin
      if (_T_6) begin
        if (io_gi_valid) begin
          if (2'h2 == jj) begin
            gamma_2_1 <= io_gi_bits_1;
          end
        end
      end
    end
    if (io_start) begin
      if (_T_6) begin
        if (io_gi_valid) begin
          if (2'h2 == jj) begin
            gamma_2_2 <= io_gi_bits_2;
          end
        end
      end
    end
    if (io_start) begin
      if (_T_6) begin
        if (io_gi_valid) begin
          if (2'h2 == jj) begin
            gamma_2_3 <= io_gi_bits_3;
          end
        end
      end
    end
    if (io_start) begin
      if (_T_6) begin
        if (io_gi_valid) begin
          if (2'h2 == jj) begin
            gamma_2_4 <= io_gi_bits_4;
          end
        end
      end
    end
    if (io_start) begin
      if (_T_6) begin
        if (io_gi_valid) begin
          if (2'h2 == jj) begin
            gamma_2_5 <= io_gi_bits_5;
          end
        end
      end
    end
    if (io_start) begin
      if (_T_6) begin
        if (io_gi_valid) begin
          if (2'h2 == jj) begin
            gamma_2_6 <= io_gi_bits_6;
          end
        end
      end
    end
    if (io_start) begin
      if (_T_6) begin
        if (io_gi_valid) begin
          if (2'h2 == jj) begin
            gamma_2_7 <= io_gi_bits_7;
          end
        end
      end
    end
    if (io_start) begin
      if (_T_6) begin
        if (io_gi_valid) begin
          if (2'h3 == jj) begin
            gamma_3_0 <= io_gi_bits_0;
          end
        end
      end
    end
    if (io_start) begin
      if (_T_6) begin
        if (io_gi_valid) begin
          if (2'h3 == jj) begin
            gamma_3_1 <= io_gi_bits_1;
          end
        end
      end
    end
    if (io_start) begin
      if (_T_6) begin
        if (io_gi_valid) begin
          if (2'h3 == jj) begin
            gamma_3_2 <= io_gi_bits_2;
          end
        end
      end
    end
    if (io_start) begin
      if (_T_6) begin
        if (io_gi_valid) begin
          if (2'h3 == jj) begin
            gamma_3_3 <= io_gi_bits_3;
          end
        end
      end
    end
    if (io_start) begin
      if (_T_6) begin
        if (io_gi_valid) begin
          if (2'h3 == jj) begin
            gamma_3_4 <= io_gi_bits_4;
          end
        end
      end
    end
    if (io_start) begin
      if (_T_6) begin
        if (io_gi_valid) begin
          if (2'h3 == jj) begin
            gamma_3_5 <= io_gi_bits_5;
          end
        end
      end
    end
    if (io_start) begin
      if (_T_6) begin
        if (io_gi_valid) begin
          if (2'h3 == jj) begin
            gamma_3_6 <= io_gi_bits_6;
          end
        end
      end
    end
    if (io_start) begin
      if (_T_6) begin
        if (io_gi_valid) begin
          if (2'h3 == jj) begin
            gamma_3_7 <= io_gi_bits_7;
          end
        end
      end
    end
    if (io_start) begin
      if (!(_T_6)) begin
        if (phase) begin
          if (_T_22) begin
            if (_T_5) begin
              if (2'h0 == _T) begin
                if (_T_5) begin
                  if (_T_57) begin
                    localWeights_0_0 <= _T_61;
                  end else begin
                    localWeights_0_0 <= _T_28;
                  end
                end else begin
                  if (2'h3 == _T) begin
                    localWeights_0_0 <= localWeights_3_0;
                  end else begin
                    if (2'h2 == _T) begin
                      localWeights_0_0 <= localWeights_2_0;
                    end else begin
                      if (2'h1 == _T) begin
                        localWeights_0_0 <= localWeights_1_0;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_start) begin
      if (!(_T_6)) begin
        if (phase) begin
          if (_T_22) begin
            if (_T_5) begin
              if (2'h0 == _T) begin
                if (_T_5) begin
                  if (_T_57) begin
                    localWeights_0_1 <= _T_65;
                  end else begin
                    localWeights_0_1 <= _T_32;
                  end
                end else begin
                  if (2'h3 == _T) begin
                    localWeights_0_1 <= localWeights_3_1;
                  end else begin
                    if (2'h2 == _T) begin
                      localWeights_0_1 <= localWeights_2_1;
                    end else begin
                      if (2'h1 == _T) begin
                        localWeights_0_1 <= localWeights_1_1;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_start) begin
      if (!(_T_6)) begin
        if (phase) begin
          if (_T_22) begin
            if (_T_5) begin
              if (2'h0 == _T) begin
                if (_T_5) begin
                  if (_T_57) begin
                    localWeights_0_2 <= _T_69;
                  end else begin
                    localWeights_0_2 <= _T_36;
                  end
                end else begin
                  if (2'h3 == _T) begin
                    localWeights_0_2 <= localWeights_3_2;
                  end else begin
                    if (2'h2 == _T) begin
                      localWeights_0_2 <= localWeights_2_2;
                    end else begin
                      if (2'h1 == _T) begin
                        localWeights_0_2 <= localWeights_1_2;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_start) begin
      if (!(_T_6)) begin
        if (phase) begin
          if (_T_22) begin
            if (_T_5) begin
              if (2'h0 == _T) begin
                if (_T_5) begin
                  if (_T_57) begin
                    localWeights_0_3 <= _T_73;
                  end else begin
                    localWeights_0_3 <= _T_40;
                  end
                end else begin
                  if (2'h3 == _T) begin
                    localWeights_0_3 <= localWeights_3_3;
                  end else begin
                    if (2'h2 == _T) begin
                      localWeights_0_3 <= localWeights_2_3;
                    end else begin
                      if (2'h1 == _T) begin
                        localWeights_0_3 <= localWeights_1_3;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_start) begin
      if (!(_T_6)) begin
        if (phase) begin
          if (_T_22) begin
            if (_T_5) begin
              if (2'h0 == _T) begin
                if (_T_5) begin
                  if (_T_57) begin
                    localWeights_0_4 <= _T_77;
                  end else begin
                    localWeights_0_4 <= _T_44;
                  end
                end else begin
                  if (2'h3 == _T) begin
                    localWeights_0_4 <= localWeights_3_4;
                  end else begin
                    if (2'h2 == _T) begin
                      localWeights_0_4 <= localWeights_2_4;
                    end else begin
                      if (2'h1 == _T) begin
                        localWeights_0_4 <= localWeights_1_4;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_start) begin
      if (!(_T_6)) begin
        if (phase) begin
          if (_T_22) begin
            if (_T_5) begin
              if (2'h0 == _T) begin
                if (_T_5) begin
                  if (_T_57) begin
                    localWeights_0_5 <= _T_81;
                  end else begin
                    localWeights_0_5 <= _T_48;
                  end
                end else begin
                  if (2'h3 == _T) begin
                    localWeights_0_5 <= localWeights_3_5;
                  end else begin
                    if (2'h2 == _T) begin
                      localWeights_0_5 <= localWeights_2_5;
                    end else begin
                      if (2'h1 == _T) begin
                        localWeights_0_5 <= localWeights_1_5;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_start) begin
      if (!(_T_6)) begin
        if (phase) begin
          if (_T_22) begin
            if (_T_5) begin
              if (2'h0 == _T) begin
                if (_T_5) begin
                  if (_T_57) begin
                    localWeights_0_6 <= _T_85;
                  end else begin
                    localWeights_0_6 <= _T_52;
                  end
                end else begin
                  if (2'h3 == _T) begin
                    localWeights_0_6 <= localWeights_3_6;
                  end else begin
                    if (2'h2 == _T) begin
                      localWeights_0_6 <= localWeights_2_6;
                    end else begin
                      if (2'h1 == _T) begin
                        localWeights_0_6 <= localWeights_1_6;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_start) begin
      if (!(_T_6)) begin
        if (phase) begin
          if (_T_22) begin
            if (_T_5) begin
              if (2'h0 == _T) begin
                if (_T_5) begin
                  if (_T_57) begin
                    localWeights_0_7 <= _T_89;
                  end else begin
                    localWeights_0_7 <= _T_56;
                  end
                end else begin
                  if (2'h3 == _T) begin
                    localWeights_0_7 <= localWeights_3_7;
                  end else begin
                    if (2'h2 == _T) begin
                      localWeights_0_7 <= localWeights_2_7;
                    end else begin
                      if (2'h1 == _T) begin
                        localWeights_0_7 <= localWeights_1_7;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_start) begin
      if (!(_T_6)) begin
        if (phase) begin
          if (_T_22) begin
            if (_T_5) begin
              if (2'h1 == _T) begin
                if (_T_5) begin
                  if (_T_57) begin
                    localWeights_1_0 <= _T_61;
                  end else begin
                    localWeights_1_0 <= _T_28;
                  end
                end else begin
                  if (2'h3 == _T) begin
                    localWeights_1_0 <= localWeights_3_0;
                  end else begin
                    if (2'h2 == _T) begin
                      localWeights_1_0 <= localWeights_2_0;
                    end else begin
                      if (!(2'h1 == _T)) begin
                        localWeights_1_0 <= localWeights_0_0;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_start) begin
      if (!(_T_6)) begin
        if (phase) begin
          if (_T_22) begin
            if (_T_5) begin
              if (2'h1 == _T) begin
                if (_T_5) begin
                  if (_T_57) begin
                    localWeights_1_1 <= _T_65;
                  end else begin
                    localWeights_1_1 <= _T_32;
                  end
                end else begin
                  if (2'h3 == _T) begin
                    localWeights_1_1 <= localWeights_3_1;
                  end else begin
                    if (2'h2 == _T) begin
                      localWeights_1_1 <= localWeights_2_1;
                    end else begin
                      if (!(2'h1 == _T)) begin
                        localWeights_1_1 <= localWeights_0_1;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_start) begin
      if (!(_T_6)) begin
        if (phase) begin
          if (_T_22) begin
            if (_T_5) begin
              if (2'h1 == _T) begin
                if (_T_5) begin
                  if (_T_57) begin
                    localWeights_1_2 <= _T_69;
                  end else begin
                    localWeights_1_2 <= _T_36;
                  end
                end else begin
                  if (2'h3 == _T) begin
                    localWeights_1_2 <= localWeights_3_2;
                  end else begin
                    if (2'h2 == _T) begin
                      localWeights_1_2 <= localWeights_2_2;
                    end else begin
                      if (!(2'h1 == _T)) begin
                        localWeights_1_2 <= localWeights_0_2;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_start) begin
      if (!(_T_6)) begin
        if (phase) begin
          if (_T_22) begin
            if (_T_5) begin
              if (2'h1 == _T) begin
                if (_T_5) begin
                  if (_T_57) begin
                    localWeights_1_3 <= _T_73;
                  end else begin
                    localWeights_1_3 <= _T_40;
                  end
                end else begin
                  if (2'h3 == _T) begin
                    localWeights_1_3 <= localWeights_3_3;
                  end else begin
                    if (2'h2 == _T) begin
                      localWeights_1_3 <= localWeights_2_3;
                    end else begin
                      if (!(2'h1 == _T)) begin
                        localWeights_1_3 <= localWeights_0_3;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_start) begin
      if (!(_T_6)) begin
        if (phase) begin
          if (_T_22) begin
            if (_T_5) begin
              if (2'h1 == _T) begin
                if (_T_5) begin
                  if (_T_57) begin
                    localWeights_1_4 <= _T_77;
                  end else begin
                    localWeights_1_4 <= _T_44;
                  end
                end else begin
                  if (2'h3 == _T) begin
                    localWeights_1_4 <= localWeights_3_4;
                  end else begin
                    if (2'h2 == _T) begin
                      localWeights_1_4 <= localWeights_2_4;
                    end else begin
                      if (!(2'h1 == _T)) begin
                        localWeights_1_4 <= localWeights_0_4;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_start) begin
      if (!(_T_6)) begin
        if (phase) begin
          if (_T_22) begin
            if (_T_5) begin
              if (2'h1 == _T) begin
                if (_T_5) begin
                  if (_T_57) begin
                    localWeights_1_5 <= _T_81;
                  end else begin
                    localWeights_1_5 <= _T_48;
                  end
                end else begin
                  if (2'h3 == _T) begin
                    localWeights_1_5 <= localWeights_3_5;
                  end else begin
                    if (2'h2 == _T) begin
                      localWeights_1_5 <= localWeights_2_5;
                    end else begin
                      if (!(2'h1 == _T)) begin
                        localWeights_1_5 <= localWeights_0_5;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_start) begin
      if (!(_T_6)) begin
        if (phase) begin
          if (_T_22) begin
            if (_T_5) begin
              if (2'h1 == _T) begin
                if (_T_5) begin
                  if (_T_57) begin
                    localWeights_1_6 <= _T_85;
                  end else begin
                    localWeights_1_6 <= _T_52;
                  end
                end else begin
                  if (2'h3 == _T) begin
                    localWeights_1_6 <= localWeights_3_6;
                  end else begin
                    if (2'h2 == _T) begin
                      localWeights_1_6 <= localWeights_2_6;
                    end else begin
                      if (!(2'h1 == _T)) begin
                        localWeights_1_6 <= localWeights_0_6;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_start) begin
      if (!(_T_6)) begin
        if (phase) begin
          if (_T_22) begin
            if (_T_5) begin
              if (2'h1 == _T) begin
                if (_T_5) begin
                  if (_T_57) begin
                    localWeights_1_7 <= _T_89;
                  end else begin
                    localWeights_1_7 <= _T_56;
                  end
                end else begin
                  if (2'h3 == _T) begin
                    localWeights_1_7 <= localWeights_3_7;
                  end else begin
                    if (2'h2 == _T) begin
                      localWeights_1_7 <= localWeights_2_7;
                    end else begin
                      if (!(2'h1 == _T)) begin
                        localWeights_1_7 <= localWeights_0_7;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_start) begin
      if (!(_T_6)) begin
        if (phase) begin
          if (_T_22) begin
            if (_T_5) begin
              if (2'h2 == _T) begin
                if (_T_5) begin
                  if (_T_57) begin
                    localWeights_2_0 <= _T_61;
                  end else begin
                    localWeights_2_0 <= _T_28;
                  end
                end else begin
                  if (2'h3 == _T) begin
                    localWeights_2_0 <= localWeights_3_0;
                  end else begin
                    if (!(2'h2 == _T)) begin
                      if (2'h1 == _T) begin
                        localWeights_2_0 <= localWeights_1_0;
                      end else begin
                        localWeights_2_0 <= localWeights_0_0;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_start) begin
      if (!(_T_6)) begin
        if (phase) begin
          if (_T_22) begin
            if (_T_5) begin
              if (2'h2 == _T) begin
                if (_T_5) begin
                  if (_T_57) begin
                    localWeights_2_1 <= _T_65;
                  end else begin
                    localWeights_2_1 <= _T_32;
                  end
                end else begin
                  if (2'h3 == _T) begin
                    localWeights_2_1 <= localWeights_3_1;
                  end else begin
                    if (!(2'h2 == _T)) begin
                      if (2'h1 == _T) begin
                        localWeights_2_1 <= localWeights_1_1;
                      end else begin
                        localWeights_2_1 <= localWeights_0_1;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_start) begin
      if (!(_T_6)) begin
        if (phase) begin
          if (_T_22) begin
            if (_T_5) begin
              if (2'h2 == _T) begin
                if (_T_5) begin
                  if (_T_57) begin
                    localWeights_2_2 <= _T_69;
                  end else begin
                    localWeights_2_2 <= _T_36;
                  end
                end else begin
                  if (2'h3 == _T) begin
                    localWeights_2_2 <= localWeights_3_2;
                  end else begin
                    if (!(2'h2 == _T)) begin
                      if (2'h1 == _T) begin
                        localWeights_2_2 <= localWeights_1_2;
                      end else begin
                        localWeights_2_2 <= localWeights_0_2;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_start) begin
      if (!(_T_6)) begin
        if (phase) begin
          if (_T_22) begin
            if (_T_5) begin
              if (2'h2 == _T) begin
                if (_T_5) begin
                  if (_T_57) begin
                    localWeights_2_3 <= _T_73;
                  end else begin
                    localWeights_2_3 <= _T_40;
                  end
                end else begin
                  if (2'h3 == _T) begin
                    localWeights_2_3 <= localWeights_3_3;
                  end else begin
                    if (!(2'h2 == _T)) begin
                      if (2'h1 == _T) begin
                        localWeights_2_3 <= localWeights_1_3;
                      end else begin
                        localWeights_2_3 <= localWeights_0_3;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_start) begin
      if (!(_T_6)) begin
        if (phase) begin
          if (_T_22) begin
            if (_T_5) begin
              if (2'h2 == _T) begin
                if (_T_5) begin
                  if (_T_57) begin
                    localWeights_2_4 <= _T_77;
                  end else begin
                    localWeights_2_4 <= _T_44;
                  end
                end else begin
                  if (2'h3 == _T) begin
                    localWeights_2_4 <= localWeights_3_4;
                  end else begin
                    if (!(2'h2 == _T)) begin
                      if (2'h1 == _T) begin
                        localWeights_2_4 <= localWeights_1_4;
                      end else begin
                        localWeights_2_4 <= localWeights_0_4;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_start) begin
      if (!(_T_6)) begin
        if (phase) begin
          if (_T_22) begin
            if (_T_5) begin
              if (2'h2 == _T) begin
                if (_T_5) begin
                  if (_T_57) begin
                    localWeights_2_5 <= _T_81;
                  end else begin
                    localWeights_2_5 <= _T_48;
                  end
                end else begin
                  if (2'h3 == _T) begin
                    localWeights_2_5 <= localWeights_3_5;
                  end else begin
                    if (!(2'h2 == _T)) begin
                      if (2'h1 == _T) begin
                        localWeights_2_5 <= localWeights_1_5;
                      end else begin
                        localWeights_2_5 <= localWeights_0_5;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_start) begin
      if (!(_T_6)) begin
        if (phase) begin
          if (_T_22) begin
            if (_T_5) begin
              if (2'h2 == _T) begin
                if (_T_5) begin
                  if (_T_57) begin
                    localWeights_2_6 <= _T_85;
                  end else begin
                    localWeights_2_6 <= _T_52;
                  end
                end else begin
                  if (2'h3 == _T) begin
                    localWeights_2_6 <= localWeights_3_6;
                  end else begin
                    if (!(2'h2 == _T)) begin
                      if (2'h1 == _T) begin
                        localWeights_2_6 <= localWeights_1_6;
                      end else begin
                        localWeights_2_6 <= localWeights_0_6;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_start) begin
      if (!(_T_6)) begin
        if (phase) begin
          if (_T_22) begin
            if (_T_5) begin
              if (2'h2 == _T) begin
                if (_T_5) begin
                  if (_T_57) begin
                    localWeights_2_7 <= _T_89;
                  end else begin
                    localWeights_2_7 <= _T_56;
                  end
                end else begin
                  if (2'h3 == _T) begin
                    localWeights_2_7 <= localWeights_3_7;
                  end else begin
                    if (!(2'h2 == _T)) begin
                      if (2'h1 == _T) begin
                        localWeights_2_7 <= localWeights_1_7;
                      end else begin
                        localWeights_2_7 <= localWeights_0_7;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_start) begin
      if (!(_T_6)) begin
        if (phase) begin
          if (_T_22) begin
            if (_T_5) begin
              if (2'h3 == _T) begin
                if (_T_5) begin
                  if (_T_57) begin
                    localWeights_3_0 <= _T_61;
                  end else begin
                    localWeights_3_0 <= _T_28;
                  end
                end else begin
                  if (!(2'h3 == _T)) begin
                    if (2'h2 == _T) begin
                      localWeights_3_0 <= localWeights_2_0;
                    end else begin
                      if (2'h1 == _T) begin
                        localWeights_3_0 <= localWeights_1_0;
                      end else begin
                        localWeights_3_0 <= localWeights_0_0;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_start) begin
      if (!(_T_6)) begin
        if (phase) begin
          if (_T_22) begin
            if (_T_5) begin
              if (2'h3 == _T) begin
                if (_T_5) begin
                  if (_T_57) begin
                    localWeights_3_1 <= _T_65;
                  end else begin
                    localWeights_3_1 <= _T_32;
                  end
                end else begin
                  if (!(2'h3 == _T)) begin
                    if (2'h2 == _T) begin
                      localWeights_3_1 <= localWeights_2_1;
                    end else begin
                      if (2'h1 == _T) begin
                        localWeights_3_1 <= localWeights_1_1;
                      end else begin
                        localWeights_3_1 <= localWeights_0_1;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_start) begin
      if (!(_T_6)) begin
        if (phase) begin
          if (_T_22) begin
            if (_T_5) begin
              if (2'h3 == _T) begin
                if (_T_5) begin
                  if (_T_57) begin
                    localWeights_3_2 <= _T_69;
                  end else begin
                    localWeights_3_2 <= _T_36;
                  end
                end else begin
                  if (!(2'h3 == _T)) begin
                    if (2'h2 == _T) begin
                      localWeights_3_2 <= localWeights_2_2;
                    end else begin
                      if (2'h1 == _T) begin
                        localWeights_3_2 <= localWeights_1_2;
                      end else begin
                        localWeights_3_2 <= localWeights_0_2;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_start) begin
      if (!(_T_6)) begin
        if (phase) begin
          if (_T_22) begin
            if (_T_5) begin
              if (2'h3 == _T) begin
                if (_T_5) begin
                  if (_T_57) begin
                    localWeights_3_3 <= _T_73;
                  end else begin
                    localWeights_3_3 <= _T_40;
                  end
                end else begin
                  if (!(2'h3 == _T)) begin
                    if (2'h2 == _T) begin
                      localWeights_3_3 <= localWeights_2_3;
                    end else begin
                      if (2'h1 == _T) begin
                        localWeights_3_3 <= localWeights_1_3;
                      end else begin
                        localWeights_3_3 <= localWeights_0_3;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_start) begin
      if (!(_T_6)) begin
        if (phase) begin
          if (_T_22) begin
            if (_T_5) begin
              if (2'h3 == _T) begin
                if (_T_5) begin
                  if (_T_57) begin
                    localWeights_3_4 <= _T_77;
                  end else begin
                    localWeights_3_4 <= _T_44;
                  end
                end else begin
                  if (!(2'h3 == _T)) begin
                    if (2'h2 == _T) begin
                      localWeights_3_4 <= localWeights_2_4;
                    end else begin
                      if (2'h1 == _T) begin
                        localWeights_3_4 <= localWeights_1_4;
                      end else begin
                        localWeights_3_4 <= localWeights_0_4;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_start) begin
      if (!(_T_6)) begin
        if (phase) begin
          if (_T_22) begin
            if (_T_5) begin
              if (2'h3 == _T) begin
                if (_T_5) begin
                  if (_T_57) begin
                    localWeights_3_5 <= _T_81;
                  end else begin
                    localWeights_3_5 <= _T_48;
                  end
                end else begin
                  if (!(2'h3 == _T)) begin
                    if (2'h2 == _T) begin
                      localWeights_3_5 <= localWeights_2_5;
                    end else begin
                      if (2'h1 == _T) begin
                        localWeights_3_5 <= localWeights_1_5;
                      end else begin
                        localWeights_3_5 <= localWeights_0_5;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_start) begin
      if (!(_T_6)) begin
        if (phase) begin
          if (_T_22) begin
            if (_T_5) begin
              if (2'h3 == _T) begin
                if (_T_5) begin
                  if (_T_57) begin
                    localWeights_3_6 <= _T_85;
                  end else begin
                    localWeights_3_6 <= _T_52;
                  end
                end else begin
                  if (!(2'h3 == _T)) begin
                    if (2'h2 == _T) begin
                      localWeights_3_6 <= localWeights_2_6;
                    end else begin
                      if (2'h1 == _T) begin
                        localWeights_3_6 <= localWeights_1_6;
                      end else begin
                        localWeights_3_6 <= localWeights_0_6;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (io_start) begin
      if (!(_T_6)) begin
        if (phase) begin
          if (_T_22) begin
            if (_T_5) begin
              if (2'h3 == _T) begin
                if (_T_5) begin
                  if (_T_57) begin
                    localWeights_3_7 <= _T_89;
                  end else begin
                    localWeights_3_7 <= _T_56;
                  end
                end else begin
                  if (!(2'h3 == _T)) begin
                    if (2'h2 == _T) begin
                      localWeights_3_7 <= localWeights_2_7;
                    end else begin
                      if (2'h1 == _T) begin
                        localWeights_3_7 <= localWeights_1_7;
                      end else begin
                        localWeights_3_7 <= localWeights_0_7;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
  end
endmodule
module Backend(
  input         clock,
  input         reset,
  input         io_start,
  output        io_done,
  output        io_res_ready,
  input         io_res_valid,
  input  [15:0] io_res_bits_0,
  input  [15:0] io_res_bits_1,
  input  [15:0] io_res_bits_2,
  input  [15:0] io_res_bits_3,
  input  [15:0] io_res_bits_4,
  input  [15:0] io_res_bits_5,
  input  [15:0] io_res_bits_6,
  input  [15:0] io_res_bits_7,
  input         io_mo_ready,
  output        io_mo_valid,
  output [15:0] io_mo_bits_bits_0,
  output [15:0] io_mo_bits_bits_1,
  output [15:0] io_mo_bits_bits_2,
  output [15:0] io_mo_bits_bits_3,
  output [15:0] io_mo_bits_bits_4,
  output [15:0] io_mo_bits_bits_5,
  output [15:0] io_mo_bits_bits_6,
  output [15:0] io_mo_bits_bits_7,
  input         io_adj_ready,
  output        io_adj_valid,
  output [15:0] io_adj_bits_0,
  output [15:0] io_adj_bits_1,
  output [15:0] io_adj_bits_2,
  output [15:0] io_adj_bits_3,
  output [15:0] io_adj_bits_4,
  output [15:0] io_adj_bits_5,
  output [15:0] io_adj_bits_6,
  output [15:0] io_adj_bits_7
);
  reg [127:0] weights [0:127]; // @[Backend.scala 32:20]
  reg [127:0] _RAND_0;
  wire [127:0] weights__T_19_data; // @[Backend.scala 32:20]
  wire [6:0] weights__T_19_addr; // @[Backend.scala 32:20]
  wire [127:0] weights__T_56_data; // @[Backend.scala 32:20]
  wire [6:0] weights__T_56_addr; // @[Backend.scala 32:20]
  wire  weights__T_56_mask; // @[Backend.scala 32:20]
  wire  weights__T_56_en; // @[Backend.scala 32:20]
  reg [1:0] _T; // @[SliceCounter.scala 7:19]
  reg [31:0] _RAND_1;
  reg [4:0] _T_1; // @[SliceCounter.scala 8:19]
  reg [31:0] _RAND_2;
  reg [4:0] _T_2; // @[SliceCounter.scala 9:19]
  reg [31:0] _RAND_3;
  reg  _T_4; // @[SliceCounter.scala 11:21]
  reg [31:0] _RAND_4;
  wire  _T_6; // @[Backend.scala 43:22]
  wire  _T_7; // @[Backend.scala 43:19]
  wire  _T_8; // @[Backend.scala 47:24]
  wire [4:0] _T_10; // @[Backend.scala 49:18]
  wire  _T_11; // @[Backend.scala 49:23]
  wire  _T_12; // @[Backend.scala 49:33]
  wire  _T_13; // @[Backend.scala 48:23]
  wire [6:0] _T_15; // @[Backend.scala 54:23]
  wire [6:0] _GEN_105; // @[Backend.scala 54:45]
  wire  _T_18; // @[Backend.scala 55:20]
  wire [127:0] _T_21;
  wire [15:0] _T_22; // @[Backend.scala 58:45]
  wire [15:0] _T_23; // @[Backend.scala 58:45]
  wire [15:0] _T_24; // @[Backend.scala 58:45]
  wire [15:0] _T_25; // @[Backend.scala 58:45]
  wire [15:0] _T_26; // @[Backend.scala 58:45]
  wire [15:0] _T_27; // @[Backend.scala 58:45]
  wire [15:0] _T_28; // @[Backend.scala 58:45]
  wire [15:0] _T_29; // @[Backend.scala 58:45]
  wire [15:0] _T_31; // @[Backend.scala 60:27]
  wire [15:0] _T_33; // @[Backend.scala 60:27]
  wire [15:0] _T_35; // @[Backend.scala 60:27]
  wire [15:0] _T_37; // @[Backend.scala 60:27]
  wire [15:0] _T_39; // @[Backend.scala 60:27]
  wire [15:0] _T_41; // @[Backend.scala 60:27]
  wire [15:0] _T_43; // @[Backend.scala 60:27]
  wire [15:0] _T_45; // @[Backend.scala 60:27]
  wire [15:0] _GEN_0; // @[Backend.scala 55:29]
  wire [15:0] _GEN_1; // @[Backend.scala 55:29]
  wire [15:0] _GEN_2; // @[Backend.scala 55:29]
  wire [15:0] _GEN_3; // @[Backend.scala 55:29]
  wire [15:0] _GEN_4; // @[Backend.scala 55:29]
  wire [15:0] _GEN_5; // @[Backend.scala 55:29]
  wire [15:0] _GEN_6; // @[Backend.scala 55:29]
  wire [15:0] _GEN_7; // @[Backend.scala 55:29]
  wire  _GEN_10; // @[Backend.scala 55:29]
  wire  _T_48; // @[Backend.scala 64:24]
  wire [63:0] _T_51; // @[Backend.scala 69:28]
  wire [63:0] _T_54; // @[Backend.scala 69:28]
  wire  _T_57; // @[SliceCounter.scala 15:9]
  wire  _T_58; // @[SliceCounter.scala 16:9]
  wire  _T_59; // @[SliceCounter.scala 15:31]
  wire  _T_60; // @[SliceCounter.scala 17:9]
  wire  _T_61; // @[SliceCounter.scala 16:22]
  wire  _T_66; // @[SliceCounter.scala 22:15]
  wire  _T_69; // @[SliceCounter.scala 26:16]
  wire  _T_72; // @[SliceCounter.scala 31:18]
  wire  _GEN_23; // @[SliceCounter.scala 31:31]
  wire  _GEN_28; // @[SliceCounter.scala 26:29]
  wire  _GEN_34; // @[SliceCounter.scala 22:37]
  wire  _GEN_66; // @[Backend.scala 49:51]
  wire  _GEN_98; // @[Backend.scala 43:32]
  wire  _T_62; // @[Backend.scala 76:28]
  wire  _T_64; // @[Backend.scala 76:13]
  wire  _T_65; // @[Backend.scala 76:13]
  wire [1:0] _T_68; // @[SliceCounter.scala 23:16]
  wire [4:0] _T_71; // @[SliceCounter.scala 27:16]
  wire [4:0] _T_74; // @[SliceCounter.scala 32:18]
  wire [4:0] _T_76; // @[SliceCounter.scala 33:18]
  wire  _GEN_38; // @[Backend.scala 49:51]
  wire  _GEN_39; // @[Backend.scala 49:51]
  wire  _GEN_106; // @[Backend.scala 76:13]
  assign weights__T_19_addr = _T_15 + _GEN_105;
  assign weights__T_19_data = weights[weights__T_19_addr]; // @[Backend.scala 32:20]
  assign weights__T_56_data = {_T_54,_T_51};
  assign weights__T_56_addr = _T_15 + _GEN_105;
  assign weights__T_56_mask = 1'h1;
  assign weights__T_56_en = _T_7 ? _T_13 : 1'h0;
  assign _T_6 = io_done == 1'h0; // @[Backend.scala 43:22]
  assign _T_7 = io_start & _T_6; // @[Backend.scala 43:19]
  assign _T_8 = io_res_valid & io_mo_ready; // @[Backend.scala 47:24]
  assign _T_10 = _T_1 - 5'h1; // @[Backend.scala 49:18]
  assign _T_11 = _T_10 != _T_2; // @[Backend.scala 49:23]
  assign _T_12 = _T_11 | io_adj_ready; // @[Backend.scala 49:33]
  assign _T_13 = _T_8 & _T_12; // @[Backend.scala 48:23]
  assign _T_15 = {_T_1, 2'h0}; // @[Backend.scala 54:23]
  assign _GEN_105 = {{5'd0}, _T}; // @[Backend.scala 54:45]
  assign _T_18 = _T_2 == 5'h0; // @[Backend.scala 55:20]
  assign _T_21 = weights__T_19_data;
  assign _T_22 = _T_21[15:0]; // @[Backend.scala 58:45]
  assign _T_23 = _T_21[31:16]; // @[Backend.scala 58:45]
  assign _T_24 = _T_21[47:32]; // @[Backend.scala 58:45]
  assign _T_25 = _T_21[63:48]; // @[Backend.scala 58:45]
  assign _T_26 = _T_21[79:64]; // @[Backend.scala 58:45]
  assign _T_27 = _T_21[95:80]; // @[Backend.scala 58:45]
  assign _T_28 = _T_21[111:96]; // @[Backend.scala 58:45]
  assign _T_29 = _T_21[127:112]; // @[Backend.scala 58:45]
  assign _T_31 = _T_22 + io_res_bits_0; // @[Backend.scala 60:27]
  assign _T_33 = _T_23 + io_res_bits_1; // @[Backend.scala 60:27]
  assign _T_35 = _T_24 + io_res_bits_2; // @[Backend.scala 60:27]
  assign _T_37 = _T_25 + io_res_bits_3; // @[Backend.scala 60:27]
  assign _T_39 = _T_26 + io_res_bits_4; // @[Backend.scala 60:27]
  assign _T_41 = _T_27 + io_res_bits_5; // @[Backend.scala 60:27]
  assign _T_43 = _T_28 + io_res_bits_6; // @[Backend.scala 60:27]
  assign _T_45 = _T_29 + io_res_bits_7; // @[Backend.scala 60:27]
  assign _GEN_0 = _T_18 ? io_res_bits_0 : _T_31; // @[Backend.scala 55:29]
  assign _GEN_1 = _T_18 ? io_res_bits_1 : _T_33; // @[Backend.scala 55:29]
  assign _GEN_2 = _T_18 ? io_res_bits_2 : _T_35; // @[Backend.scala 55:29]
  assign _GEN_3 = _T_18 ? io_res_bits_3 : _T_37; // @[Backend.scala 55:29]
  assign _GEN_4 = _T_18 ? io_res_bits_4 : _T_39; // @[Backend.scala 55:29]
  assign _GEN_5 = _T_18 ? io_res_bits_5 : _T_41; // @[Backend.scala 55:29]
  assign _GEN_6 = _T_18 ? io_res_bits_6 : _T_43; // @[Backend.scala 55:29]
  assign _GEN_7 = _T_18 ? io_res_bits_7 : _T_45; // @[Backend.scala 55:29]
  assign _GEN_10 = _T_18 ? 1'h0 : 1'h1; // @[Backend.scala 55:29]
  assign _T_48 = _T_10 == _T_2; // @[Backend.scala 64:24]
  assign _T_51 = {_GEN_3,_GEN_2,_GEN_1,_GEN_0}; // @[Backend.scala 69:28]
  assign _T_54 = {_GEN_7,_GEN_6,_GEN_5,_GEN_4}; // @[Backend.scala 69:28]
  assign _T_57 = _T == 2'h2; // @[SliceCounter.scala 15:9]
  assign _T_58 = _T_1 == 5'h17; // @[SliceCounter.scala 16:9]
  assign _T_59 = _T_57 & _T_58; // @[SliceCounter.scala 15:31]
  assign _T_60 = _T_2 == 5'h16; // @[SliceCounter.scala 17:9]
  assign _T_61 = _T_59 & _T_60; // @[SliceCounter.scala 16:22]
  assign _T_66 = _T != 2'h2; // @[SliceCounter.scala 22:15]
  assign _T_69 = _T_1 != 5'h17; // @[SliceCounter.scala 26:16]
  assign _T_72 = _T_2 != 5'h16; // @[SliceCounter.scala 31:18]
  assign _GEN_23 = _T_72 ? 1'h0 : 1'h1; // @[SliceCounter.scala 31:31]
  assign _GEN_28 = _T_69 ? 1'h0 : _GEN_23; // @[SliceCounter.scala 26:29]
  assign _GEN_34 = _T_66 ? 1'h0 : _GEN_28; // @[SliceCounter.scala 22:37]
  assign _GEN_66 = _T_13 ? _GEN_34 : 1'h0; // @[Backend.scala 49:51]
  assign _GEN_98 = _T_7 ? _GEN_66 : 1'h0; // @[Backend.scala 43:32]
  assign _T_62 = _GEN_98 == _T_61; // @[Backend.scala 76:28]
  assign _T_64 = _T_62 | reset; // @[Backend.scala 76:13]
  assign _T_65 = _T_64 == 1'h0; // @[Backend.scala 76:13]
  assign _T_68 = _T + 2'h1; // @[SliceCounter.scala 23:16]
  assign _T_71 = _T_1 + 5'h1; // @[SliceCounter.scala 27:16]
  assign _T_74 = _T_2 + 5'h1; // @[SliceCounter.scala 32:18]
  assign _T_76 = _T_2 + 5'h2; // @[SliceCounter.scala 33:18]
  assign _GEN_38 = _T_13 ? _GEN_10 : 1'h0; // @[Backend.scala 49:51]
  assign _GEN_39 = _T_13 ? _T_48 : 1'h0; // @[Backend.scala 49:51]
  assign io_done = _T_4; // @[Backend.scala 34:11]
  assign io_res_ready = _T_7 ? _T_13 : 1'h0; // @[Decoupled.scala 69:20 Backend.scala 50:20]
  assign io_mo_valid = _T_7 ? _T_13 : 1'h0; // @[Decoupled.scala 53:20 Backend.scala 71:19]
  assign io_mo_bits_bits_0 = io_res_bits_0; // @[Backend.scala 73:23]
  assign io_mo_bits_bits_1 = io_res_bits_1; // @[Backend.scala 73:23]
  assign io_mo_bits_bits_2 = io_res_bits_2; // @[Backend.scala 73:23]
  assign io_mo_bits_bits_3 = io_res_bits_3; // @[Backend.scala 73:23]
  assign io_mo_bits_bits_4 = io_res_bits_4; // @[Backend.scala 73:23]
  assign io_mo_bits_bits_5 = io_res_bits_5; // @[Backend.scala 73:23]
  assign io_mo_bits_bits_6 = io_res_bits_6; // @[Backend.scala 73:23]
  assign io_mo_bits_bits_7 = io_res_bits_7; // @[Backend.scala 73:23]
  assign io_adj_valid = _T_7 ? _GEN_39 : 1'h0; // @[Decoupled.scala 53:20 Backend.scala 65:22]
  assign io_adj_bits_0 = _T_18 ? io_res_bits_0 : _T_31; // @[Backend.scala 66:21]
  assign io_adj_bits_1 = _T_18 ? io_res_bits_1 : _T_33; // @[Backend.scala 66:21]
  assign io_adj_bits_2 = _T_18 ? io_res_bits_2 : _T_35; // @[Backend.scala 66:21]
  assign io_adj_bits_3 = _T_18 ? io_res_bits_3 : _T_37; // @[Backend.scala 66:21]
  assign io_adj_bits_4 = _T_18 ? io_res_bits_4 : _T_39; // @[Backend.scala 66:21]
  assign io_adj_bits_5 = _T_18 ? io_res_bits_5 : _T_41; // @[Backend.scala 66:21]
  assign io_adj_bits_6 = _T_18 ? io_res_bits_6 : _T_43; // @[Backend.scala 66:21]
  assign io_adj_bits_7 = _T_18 ? io_res_bits_7 : _T_45; // @[Backend.scala 66:21]
  assign _GEN_106 = _T_7 & _T_13; // @[Backend.scala 76:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {4{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    weights[initvar] = _RAND_0[127:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_1 = _RAND_2[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_2 = _RAND_3[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_4 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(weights__T_56_en & weights__T_56_mask) begin
      weights[weights__T_56_addr] <= weights__T_56_data; // @[Backend.scala 32:20]
    end
    if (reset) begin
      _T <= 2'h0;
    end else begin
      if (_T_7) begin
        if (_T_13) begin
          if (_T_66) begin
            _T <= _T_68;
          end else begin
            _T <= 2'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_1 <= 5'h1;
    end else begin
      if (_T_7) begin
        if (_T_13) begin
          if (!(_T_66)) begin
            if (_T_69) begin
              _T_1 <= _T_71;
            end else begin
              if (_T_72) begin
                _T_1 <= _T_76;
              end else begin
                _T_1 <= 5'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_2 <= 5'h0;
    end else begin
      if (_T_7) begin
        if (_T_13) begin
          if (!(_T_66)) begin
            if (!(_T_69)) begin
              if (_T_72) begin
                _T_2 <= _T_74;
              end else begin
                _T_2 <= 5'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_4 <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_13) begin
          if (!(_T_66)) begin
            if (!(_T_69)) begin
              if (!(_T_72)) begin
                _T_4 <= 1'h1;
              end
            end
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_106 & _T_65) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Backend.scala:76 assert( sc2.doneWire === sc2.lastMessage)\n"); // @[Backend.scala 76:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_106 & _T_65) begin
          $fatal; // @[Backend.scala 76:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Accumulator(
  input         clock,
  input         reset,
  output        io_mi0_ready,
  input         io_mi0_valid,
  input  [15:0] io_mi0_bits_0,
  input  [15:0] io_mi0_bits_1,
  input  [15:0] io_mi0_bits_2,
  input  [15:0] io_mi0_bits_3,
  input  [15:0] io_mi0_bits_4,
  input  [15:0] io_mi0_bits_5,
  input  [15:0] io_mi0_bits_6,
  input  [15:0] io_mi0_bits_7,
  input         io_a0_ready,
  output        io_a0_valid,
  output [15:0] io_a0_bits_0,
  output [15:0] io_a0_bits_1,
  output [15:0] io_a0_bits_2,
  output [15:0] io_a0_bits_3,
  output [15:0] io_a0_bits_4,
  output [15:0] io_a0_bits_5,
  output [15:0] io_a0_bits_6,
  output [15:0] io_a0_bits_7
);
  reg [1:0] _T; // @[SliceCounter.scala 7:19]
  reg [31:0] _RAND_0;
  reg [4:0] _T_1; // @[SliceCounter.scala 8:19]
  reg [31:0] _RAND_1;
  reg [4:0] _T_2; // @[SliceCounter.scala 9:19]
  reg [31:0] _RAND_2;
  reg  _T_5; // @[SliceCounter.scala 12:24]
  reg [31:0] _RAND_3;
  reg [15:0] localWeights_0_0; // @[Accumulator.scala 16:25]
  reg [31:0] _RAND_4;
  reg [15:0] localWeights_0_1; // @[Accumulator.scala 16:25]
  reg [31:0] _RAND_5;
  reg [15:0] localWeights_0_2; // @[Accumulator.scala 16:25]
  reg [31:0] _RAND_6;
  reg [15:0] localWeights_0_3; // @[Accumulator.scala 16:25]
  reg [31:0] _RAND_7;
  reg [15:0] localWeights_0_4; // @[Accumulator.scala 16:25]
  reg [31:0] _RAND_8;
  reg [15:0] localWeights_0_5; // @[Accumulator.scala 16:25]
  reg [31:0] _RAND_9;
  reg [15:0] localWeights_0_6; // @[Accumulator.scala 16:25]
  reg [31:0] _RAND_10;
  reg [15:0] localWeights_0_7; // @[Accumulator.scala 16:25]
  reg [31:0] _RAND_11;
  reg [15:0] localWeights_1_0; // @[Accumulator.scala 16:25]
  reg [31:0] _RAND_12;
  reg [15:0] localWeights_1_1; // @[Accumulator.scala 16:25]
  reg [31:0] _RAND_13;
  reg [15:0] localWeights_1_2; // @[Accumulator.scala 16:25]
  reg [31:0] _RAND_14;
  reg [15:0] localWeights_1_3; // @[Accumulator.scala 16:25]
  reg [31:0] _RAND_15;
  reg [15:0] localWeights_1_4; // @[Accumulator.scala 16:25]
  reg [31:0] _RAND_16;
  reg [15:0] localWeights_1_5; // @[Accumulator.scala 16:25]
  reg [31:0] _RAND_17;
  reg [15:0] localWeights_1_6; // @[Accumulator.scala 16:25]
  reg [31:0] _RAND_18;
  reg [15:0] localWeights_1_7; // @[Accumulator.scala 16:25]
  reg [31:0] _RAND_19;
  reg [15:0] localWeights_2_0; // @[Accumulator.scala 16:25]
  reg [31:0] _RAND_20;
  reg [15:0] localWeights_2_1; // @[Accumulator.scala 16:25]
  reg [31:0] _RAND_21;
  reg [15:0] localWeights_2_2; // @[Accumulator.scala 16:25]
  reg [31:0] _RAND_22;
  reg [15:0] localWeights_2_3; // @[Accumulator.scala 16:25]
  reg [31:0] _RAND_23;
  reg [15:0] localWeights_2_4; // @[Accumulator.scala 16:25]
  reg [31:0] _RAND_24;
  reg [15:0] localWeights_2_5; // @[Accumulator.scala 16:25]
  reg [31:0] _RAND_25;
  reg [15:0] localWeights_2_6; // @[Accumulator.scala 16:25]
  reg [31:0] _RAND_26;
  reg [15:0] localWeights_2_7; // @[Accumulator.scala 16:25]
  reg [31:0] _RAND_27;
  reg [15:0] localWeights_3_0; // @[Accumulator.scala 16:25]
  reg [31:0] _RAND_28;
  reg [15:0] localWeights_3_1; // @[Accumulator.scala 16:25]
  reg [31:0] _RAND_29;
  reg [15:0] localWeights_3_2; // @[Accumulator.scala 16:25]
  reg [31:0] _RAND_30;
  reg [15:0] localWeights_3_3; // @[Accumulator.scala 16:25]
  reg [31:0] _RAND_31;
  reg [15:0] localWeights_3_4; // @[Accumulator.scala 16:25]
  reg [31:0] _RAND_32;
  reg [15:0] localWeights_3_5; // @[Accumulator.scala 16:25]
  reg [31:0] _RAND_33;
  reg [15:0] localWeights_3_6; // @[Accumulator.scala 16:25]
  reg [31:0] _RAND_34;
  reg [15:0] localWeights_3_7; // @[Accumulator.scala 16:25]
  reg [31:0] _RAND_35;
  wire  _T_6; // @[Accumulator.scala 22:48]
  wire  _T_7; // @[Accumulator.scala 22:39]
  wire  _T_8; // @[Accumulator.scala 22:23]
  wire [15:0] _GEN_8; // @[Accumulator.scala 28:49]
  wire [15:0] _GEN_9; // @[Accumulator.scala 28:49]
  wire [15:0] _GEN_10; // @[Accumulator.scala 28:49]
  wire [15:0] _GEN_11; // @[Accumulator.scala 28:49]
  wire [15:0] _GEN_12; // @[Accumulator.scala 28:49]
  wire [15:0] _GEN_13; // @[Accumulator.scala 28:49]
  wire [15:0] _GEN_14; // @[Accumulator.scala 28:49]
  wire [15:0] _GEN_15; // @[Accumulator.scala 28:49]
  wire [15:0] _GEN_16; // @[Accumulator.scala 28:49]
  wire [15:0] _GEN_17; // @[Accumulator.scala 28:49]
  wire [15:0] _GEN_18; // @[Accumulator.scala 28:49]
  wire [15:0] _GEN_19; // @[Accumulator.scala 28:49]
  wire [15:0] _GEN_20; // @[Accumulator.scala 28:49]
  wire [15:0] _GEN_21; // @[Accumulator.scala 28:49]
  wire [15:0] _GEN_22; // @[Accumulator.scala 28:49]
  wire [15:0] _GEN_23; // @[Accumulator.scala 28:49]
  wire [15:0] _GEN_24; // @[Accumulator.scala 28:49]
  wire [15:0] _GEN_25; // @[Accumulator.scala 28:49]
  wire [15:0] _GEN_26; // @[Accumulator.scala 28:49]
  wire [15:0] _GEN_27; // @[Accumulator.scala 28:49]
  wire [15:0] _GEN_28; // @[Accumulator.scala 28:49]
  wire [15:0] _GEN_29; // @[Accumulator.scala 28:49]
  wire [15:0] _GEN_30; // @[Accumulator.scala 28:49]
  wire [15:0] _GEN_31; // @[Accumulator.scala 28:49]
  wire [15:0] _T_10; // @[Accumulator.scala 28:49]
  wire [15:0] _T_12; // @[Accumulator.scala 28:49]
  wire [15:0] _T_14; // @[Accumulator.scala 28:49]
  wire [15:0] _T_16; // @[Accumulator.scala 28:49]
  wire [15:0] _T_18; // @[Accumulator.scala 28:49]
  wire [15:0] _T_20; // @[Accumulator.scala 28:49]
  wire [15:0] _T_22; // @[Accumulator.scala 28:49]
  wire [15:0] _T_24; // @[Accumulator.scala 28:49]
  wire  _T_25; // @[Accumulator.scala 32:18]
  wire  _T_26; // @[SliceCounter.scala 22:15]
  wire [1:0] _T_28; // @[SliceCounter.scala 23:16]
  wire [4:0] _T_31; // @[SliceCounter.scala 27:16]
  wire  _T_32; // @[SliceCounter.scala 31:18]
  wire [4:0] _T_34; // @[SliceCounter.scala 32:18]
  wire [4:0] _T_36; // @[SliceCounter.scala 33:18]
  assign _T_6 = _T_1 != 5'h17; // @[Accumulator.scala 22:48]
  assign _T_7 = io_a0_ready | _T_6; // @[Accumulator.scala 22:39]
  assign _T_8 = io_mi0_valid & _T_7; // @[Accumulator.scala 22:23]
  assign _GEN_8 = 2'h1 == _T ? localWeights_1_0 : localWeights_0_0; // @[Accumulator.scala 28:49]
  assign _GEN_9 = 2'h1 == _T ? localWeights_1_1 : localWeights_0_1; // @[Accumulator.scala 28:49]
  assign _GEN_10 = 2'h1 == _T ? localWeights_1_2 : localWeights_0_2; // @[Accumulator.scala 28:49]
  assign _GEN_11 = 2'h1 == _T ? localWeights_1_3 : localWeights_0_3; // @[Accumulator.scala 28:49]
  assign _GEN_12 = 2'h1 == _T ? localWeights_1_4 : localWeights_0_4; // @[Accumulator.scala 28:49]
  assign _GEN_13 = 2'h1 == _T ? localWeights_1_5 : localWeights_0_5; // @[Accumulator.scala 28:49]
  assign _GEN_14 = 2'h1 == _T ? localWeights_1_6 : localWeights_0_6; // @[Accumulator.scala 28:49]
  assign _GEN_15 = 2'h1 == _T ? localWeights_1_7 : localWeights_0_7; // @[Accumulator.scala 28:49]
  assign _GEN_16 = 2'h2 == _T ? localWeights_2_0 : _GEN_8; // @[Accumulator.scala 28:49]
  assign _GEN_17 = 2'h2 == _T ? localWeights_2_1 : _GEN_9; // @[Accumulator.scala 28:49]
  assign _GEN_18 = 2'h2 == _T ? localWeights_2_2 : _GEN_10; // @[Accumulator.scala 28:49]
  assign _GEN_19 = 2'h2 == _T ? localWeights_2_3 : _GEN_11; // @[Accumulator.scala 28:49]
  assign _GEN_20 = 2'h2 == _T ? localWeights_2_4 : _GEN_12; // @[Accumulator.scala 28:49]
  assign _GEN_21 = 2'h2 == _T ? localWeights_2_5 : _GEN_13; // @[Accumulator.scala 28:49]
  assign _GEN_22 = 2'h2 == _T ? localWeights_2_6 : _GEN_14; // @[Accumulator.scala 28:49]
  assign _GEN_23 = 2'h2 == _T ? localWeights_2_7 : _GEN_15; // @[Accumulator.scala 28:49]
  assign _GEN_24 = 2'h3 == _T ? localWeights_3_0 : _GEN_16; // @[Accumulator.scala 28:49]
  assign _GEN_25 = 2'h3 == _T ? localWeights_3_1 : _GEN_17; // @[Accumulator.scala 28:49]
  assign _GEN_26 = 2'h3 == _T ? localWeights_3_2 : _GEN_18; // @[Accumulator.scala 28:49]
  assign _GEN_27 = 2'h3 == _T ? localWeights_3_3 : _GEN_19; // @[Accumulator.scala 28:49]
  assign _GEN_28 = 2'h3 == _T ? localWeights_3_4 : _GEN_20; // @[Accumulator.scala 28:49]
  assign _GEN_29 = 2'h3 == _T ? localWeights_3_5 : _GEN_21; // @[Accumulator.scala 28:49]
  assign _GEN_30 = 2'h3 == _T ? localWeights_3_6 : _GEN_22; // @[Accumulator.scala 28:49]
  assign _GEN_31 = 2'h3 == _T ? localWeights_3_7 : _GEN_23; // @[Accumulator.scala 28:49]
  assign _T_10 = _GEN_24 + io_mi0_bits_0; // @[Accumulator.scala 28:49]
  assign _T_12 = _GEN_25 + io_mi0_bits_1; // @[Accumulator.scala 28:49]
  assign _T_14 = _GEN_26 + io_mi0_bits_2; // @[Accumulator.scala 28:49]
  assign _T_16 = _GEN_27 + io_mi0_bits_3; // @[Accumulator.scala 28:49]
  assign _T_18 = _GEN_28 + io_mi0_bits_4; // @[Accumulator.scala 28:49]
  assign _T_20 = _GEN_29 + io_mi0_bits_5; // @[Accumulator.scala 28:49]
  assign _T_22 = _GEN_30 + io_mi0_bits_6; // @[Accumulator.scala 28:49]
  assign _T_24 = _GEN_31 + io_mi0_bits_7; // @[Accumulator.scala 28:49]
  assign _T_25 = _T_1 == 5'h17; // @[Accumulator.scala 32:18]
  assign _T_26 = _T != 2'h2; // @[SliceCounter.scala 22:15]
  assign _T_28 = _T + 2'h1; // @[SliceCounter.scala 23:16]
  assign _T_31 = _T_1 + 5'h1; // @[SliceCounter.scala 27:16]
  assign _T_32 = _T_2 != 5'h16; // @[SliceCounter.scala 31:18]
  assign _T_34 = _T_2 + 5'h1; // @[SliceCounter.scala 32:18]
  assign _T_36 = _T_2 + 5'h2; // @[SliceCounter.scala 33:18]
  assign io_mi0_ready = io_mi0_valid & _T_7; // @[Decoupled.scala 69:20 Accumulator.scala 23:18]
  assign io_a0_valid = _T_8 ? _T_25 : 1'h0; // @[Decoupled.scala 53:20 Accumulator.scala 33:19]
  assign io_a0_bits_0 = _T_5 ? io_mi0_bits_0 : _T_10; // @[Accumulator.scala 34:18]
  assign io_a0_bits_1 = _T_5 ? io_mi0_bits_1 : _T_12; // @[Accumulator.scala 34:18]
  assign io_a0_bits_2 = _T_5 ? io_mi0_bits_2 : _T_14; // @[Accumulator.scala 34:18]
  assign io_a0_bits_3 = _T_5 ? io_mi0_bits_3 : _T_16; // @[Accumulator.scala 34:18]
  assign io_a0_bits_4 = _T_5 ? io_mi0_bits_4 : _T_18; // @[Accumulator.scala 34:18]
  assign io_a0_bits_5 = _T_5 ? io_mi0_bits_5 : _T_20; // @[Accumulator.scala 34:18]
  assign io_a0_bits_6 = _T_5 ? io_mi0_bits_6 : _T_22; // @[Accumulator.scala 34:18]
  assign io_a0_bits_7 = _T_5 ? io_mi0_bits_7 : _T_24; // @[Accumulator.scala 34:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1 = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_2 = _RAND_2[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_5 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  localWeights_0_0 = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  localWeights_0_1 = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  localWeights_0_2 = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  localWeights_0_3 = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  localWeights_0_4 = _RAND_8[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  localWeights_0_5 = _RAND_9[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  localWeights_0_6 = _RAND_10[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  localWeights_0_7 = _RAND_11[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  localWeights_1_0 = _RAND_12[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  localWeights_1_1 = _RAND_13[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  localWeights_1_2 = _RAND_14[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  localWeights_1_3 = _RAND_15[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  localWeights_1_4 = _RAND_16[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  localWeights_1_5 = _RAND_17[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  localWeights_1_6 = _RAND_18[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  localWeights_1_7 = _RAND_19[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  localWeights_2_0 = _RAND_20[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  localWeights_2_1 = _RAND_21[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  localWeights_2_2 = _RAND_22[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  localWeights_2_3 = _RAND_23[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  localWeights_2_4 = _RAND_24[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  localWeights_2_5 = _RAND_25[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  localWeights_2_6 = _RAND_26[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  localWeights_2_7 = _RAND_27[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  localWeights_3_0 = _RAND_28[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  localWeights_3_1 = _RAND_29[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  localWeights_3_2 = _RAND_30[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  localWeights_3_3 = _RAND_31[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  localWeights_3_4 = _RAND_32[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  localWeights_3_5 = _RAND_33[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  localWeights_3_6 = _RAND_34[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  localWeights_3_7 = _RAND_35[15:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T <= 2'h0;
    end else begin
      if (_T_8) begin
        if (_T_26) begin
          _T <= _T_28;
        end else begin
          _T <= 2'h0;
        end
      end
    end
    if (reset) begin
      _T_1 <= 5'h1;
    end else begin
      if (_T_8) begin
        if (!(_T_26)) begin
          if (_T_6) begin
            _T_1 <= _T_31;
          end else begin
            if (_T_32) begin
              _T_1 <= _T_36;
            end else begin
              _T_1 <= 5'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      _T_2 <= 5'h0;
    end else begin
      if (_T_8) begin
        if (!(_T_26)) begin
          if (!(_T_6)) begin
            if (_T_32) begin
              _T_2 <= _T_34;
            end else begin
              _T_2 <= 5'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      _T_5 <= 1'h1;
    end else begin
      if (_T_8) begin
        if (!(_T_26)) begin
          if (_T_6) begin
            _T_5 <= 1'h0;
          end else begin
            _T_5 <= 1'h1;
          end
        end
      end
    end
    if (_T_8) begin
      if (!(_T_25)) begin
        if (2'h0 == _T) begin
          if (_T_5) begin
            localWeights_0_0 <= io_mi0_bits_0;
          end else begin
            localWeights_0_0 <= _T_10;
          end
        end
      end
    end
    if (_T_8) begin
      if (!(_T_25)) begin
        if (2'h0 == _T) begin
          if (_T_5) begin
            localWeights_0_1 <= io_mi0_bits_1;
          end else begin
            localWeights_0_1 <= _T_12;
          end
        end
      end
    end
    if (_T_8) begin
      if (!(_T_25)) begin
        if (2'h0 == _T) begin
          if (_T_5) begin
            localWeights_0_2 <= io_mi0_bits_2;
          end else begin
            localWeights_0_2 <= _T_14;
          end
        end
      end
    end
    if (_T_8) begin
      if (!(_T_25)) begin
        if (2'h0 == _T) begin
          if (_T_5) begin
            localWeights_0_3 <= io_mi0_bits_3;
          end else begin
            localWeights_0_3 <= _T_16;
          end
        end
      end
    end
    if (_T_8) begin
      if (!(_T_25)) begin
        if (2'h0 == _T) begin
          if (_T_5) begin
            localWeights_0_4 <= io_mi0_bits_4;
          end else begin
            localWeights_0_4 <= _T_18;
          end
        end
      end
    end
    if (_T_8) begin
      if (!(_T_25)) begin
        if (2'h0 == _T) begin
          if (_T_5) begin
            localWeights_0_5 <= io_mi0_bits_5;
          end else begin
            localWeights_0_5 <= _T_20;
          end
        end
      end
    end
    if (_T_8) begin
      if (!(_T_25)) begin
        if (2'h0 == _T) begin
          if (_T_5) begin
            localWeights_0_6 <= io_mi0_bits_6;
          end else begin
            localWeights_0_6 <= _T_22;
          end
        end
      end
    end
    if (_T_8) begin
      if (!(_T_25)) begin
        if (2'h0 == _T) begin
          if (_T_5) begin
            localWeights_0_7 <= io_mi0_bits_7;
          end else begin
            localWeights_0_7 <= _T_24;
          end
        end
      end
    end
    if (_T_8) begin
      if (!(_T_25)) begin
        if (2'h1 == _T) begin
          if (_T_5) begin
            localWeights_1_0 <= io_mi0_bits_0;
          end else begin
            localWeights_1_0 <= _T_10;
          end
        end
      end
    end
    if (_T_8) begin
      if (!(_T_25)) begin
        if (2'h1 == _T) begin
          if (_T_5) begin
            localWeights_1_1 <= io_mi0_bits_1;
          end else begin
            localWeights_1_1 <= _T_12;
          end
        end
      end
    end
    if (_T_8) begin
      if (!(_T_25)) begin
        if (2'h1 == _T) begin
          if (_T_5) begin
            localWeights_1_2 <= io_mi0_bits_2;
          end else begin
            localWeights_1_2 <= _T_14;
          end
        end
      end
    end
    if (_T_8) begin
      if (!(_T_25)) begin
        if (2'h1 == _T) begin
          if (_T_5) begin
            localWeights_1_3 <= io_mi0_bits_3;
          end else begin
            localWeights_1_3 <= _T_16;
          end
        end
      end
    end
    if (_T_8) begin
      if (!(_T_25)) begin
        if (2'h1 == _T) begin
          if (_T_5) begin
            localWeights_1_4 <= io_mi0_bits_4;
          end else begin
            localWeights_1_4 <= _T_18;
          end
        end
      end
    end
    if (_T_8) begin
      if (!(_T_25)) begin
        if (2'h1 == _T) begin
          if (_T_5) begin
            localWeights_1_5 <= io_mi0_bits_5;
          end else begin
            localWeights_1_5 <= _T_20;
          end
        end
      end
    end
    if (_T_8) begin
      if (!(_T_25)) begin
        if (2'h1 == _T) begin
          if (_T_5) begin
            localWeights_1_6 <= io_mi0_bits_6;
          end else begin
            localWeights_1_6 <= _T_22;
          end
        end
      end
    end
    if (_T_8) begin
      if (!(_T_25)) begin
        if (2'h1 == _T) begin
          if (_T_5) begin
            localWeights_1_7 <= io_mi0_bits_7;
          end else begin
            localWeights_1_7 <= _T_24;
          end
        end
      end
    end
    if (_T_8) begin
      if (!(_T_25)) begin
        if (2'h2 == _T) begin
          if (_T_5) begin
            localWeights_2_0 <= io_mi0_bits_0;
          end else begin
            localWeights_2_0 <= _T_10;
          end
        end
      end
    end
    if (_T_8) begin
      if (!(_T_25)) begin
        if (2'h2 == _T) begin
          if (_T_5) begin
            localWeights_2_1 <= io_mi0_bits_1;
          end else begin
            localWeights_2_1 <= _T_12;
          end
        end
      end
    end
    if (_T_8) begin
      if (!(_T_25)) begin
        if (2'h2 == _T) begin
          if (_T_5) begin
            localWeights_2_2 <= io_mi0_bits_2;
          end else begin
            localWeights_2_2 <= _T_14;
          end
        end
      end
    end
    if (_T_8) begin
      if (!(_T_25)) begin
        if (2'h2 == _T) begin
          if (_T_5) begin
            localWeights_2_3 <= io_mi0_bits_3;
          end else begin
            localWeights_2_3 <= _T_16;
          end
        end
      end
    end
    if (_T_8) begin
      if (!(_T_25)) begin
        if (2'h2 == _T) begin
          if (_T_5) begin
            localWeights_2_4 <= io_mi0_bits_4;
          end else begin
            localWeights_2_4 <= _T_18;
          end
        end
      end
    end
    if (_T_8) begin
      if (!(_T_25)) begin
        if (2'h2 == _T) begin
          if (_T_5) begin
            localWeights_2_5 <= io_mi0_bits_5;
          end else begin
            localWeights_2_5 <= _T_20;
          end
        end
      end
    end
    if (_T_8) begin
      if (!(_T_25)) begin
        if (2'h2 == _T) begin
          if (_T_5) begin
            localWeights_2_6 <= io_mi0_bits_6;
          end else begin
            localWeights_2_6 <= _T_22;
          end
        end
      end
    end
    if (_T_8) begin
      if (!(_T_25)) begin
        if (2'h2 == _T) begin
          if (_T_5) begin
            localWeights_2_7 <= io_mi0_bits_7;
          end else begin
            localWeights_2_7 <= _T_24;
          end
        end
      end
    end
    if (_T_8) begin
      if (!(_T_25)) begin
        if (2'h3 == _T) begin
          if (_T_5) begin
            localWeights_3_0 <= io_mi0_bits_0;
          end else begin
            localWeights_3_0 <= _T_10;
          end
        end
      end
    end
    if (_T_8) begin
      if (!(_T_25)) begin
        if (2'h3 == _T) begin
          if (_T_5) begin
            localWeights_3_1 <= io_mi0_bits_1;
          end else begin
            localWeights_3_1 <= _T_12;
          end
        end
      end
    end
    if (_T_8) begin
      if (!(_T_25)) begin
        if (2'h3 == _T) begin
          if (_T_5) begin
            localWeights_3_2 <= io_mi0_bits_2;
          end else begin
            localWeights_3_2 <= _T_14;
          end
        end
      end
    end
    if (_T_8) begin
      if (!(_T_25)) begin
        if (2'h3 == _T) begin
          if (_T_5) begin
            localWeights_3_3 <= io_mi0_bits_3;
          end else begin
            localWeights_3_3 <= _T_16;
          end
        end
      end
    end
    if (_T_8) begin
      if (!(_T_25)) begin
        if (2'h3 == _T) begin
          if (_T_5) begin
            localWeights_3_4 <= io_mi0_bits_4;
          end else begin
            localWeights_3_4 <= _T_18;
          end
        end
      end
    end
    if (_T_8) begin
      if (!(_T_25)) begin
        if (2'h3 == _T) begin
          if (_T_5) begin
            localWeights_3_5 <= io_mi0_bits_5;
          end else begin
            localWeights_3_5 <= _T_20;
          end
        end
      end
    end
    if (_T_8) begin
      if (!(_T_25)) begin
        if (2'h3 == _T) begin
          if (_T_5) begin
            localWeights_3_6 <= io_mi0_bits_6;
          end else begin
            localWeights_3_6 <= _T_22;
          end
        end
      end
    end
    if (_T_8) begin
      if (!(_T_25)) begin
        if (2'h3 == _T) begin
          if (_T_5) begin
            localWeights_3_7 <= io_mi0_bits_7;
          end else begin
            localWeights_3_7 <= _T_24;
          end
        end
      end
    end
  end
endmodule
module MAC(
  input         clock,
  input         io_en,
  input  [15:0] io_a,
  input  [15:0] io_b,
  input  [31:0] io_o,
  output [31:0] io_r
);
  reg [15:0] a2; // @[loaf.scala 72:15]
  reg [31:0] _RAND_0;
  reg [15:0] a3; // @[loaf.scala 73:15]
  reg [31:0] _RAND_1;
  reg [15:0] a4; // @[loaf.scala 74:15]
  reg [31:0] _RAND_2;
  reg [15:0] b2; // @[loaf.scala 75:15]
  reg [31:0] _RAND_3;
  reg [15:0] b3; // @[loaf.scala 76:15]
  reg [31:0] _RAND_4;
  reg [15:0] b4; // @[loaf.scala 77:15]
  reg [31:0] _RAND_5;
  reg [31:0] o2; // @[loaf.scala 78:15]
  reg [31:0] _RAND_6;
  reg [31:0] o3; // @[loaf.scala 79:15]
  reg [31:0] _RAND_7;
  reg [31:0] o4; // @[loaf.scala 80:15]
  reg [31:0] _RAND_8;
  reg [31:0] r5; // @[loaf.scala 82:15]
  reg [31:0] _RAND_9;
  reg [31:0] r6; // @[loaf.scala 83:15]
  reg [31:0] _RAND_10;
  wire [31:0] _T; // @[loaf.scala 95:15]
  wire [31:0] _T_1; // @[loaf.scala 95:21]
  wire [31:0] _T_3; // @[loaf.scala 95:28]
  wire [31:0] _T_4; // @[loaf.scala 95:28]
  assign _T = a4 * b4; // @[loaf.scala 95:15]
  assign _T_1 = $signed(_T); // @[loaf.scala 95:21]
  assign _T_3 = $signed(_T_1) + $signed(o4); // @[loaf.scala 95:28]
  assign _T_4 = $signed(_T_3); // @[loaf.scala 95:28]
  assign io_r = r6; // @[loaf.scala 99:8]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  a2 = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  a3 = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  a4 = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  b2 = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  b3 = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  b4 = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  o2 = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  o3 = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  o4 = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  r5 = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  r6 = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (io_en) begin
      a2 <= io_a;
    end
    if (io_en) begin
      a3 <= a2;
    end
    if (io_en) begin
      a4 <= a3;
    end
    if (io_en) begin
      b2 <= io_b;
    end
    if (io_en) begin
      b3 <= b2;
    end
    if (io_en) begin
      b4 <= b3;
    end
    if (io_en) begin
      o2 <= io_o;
    end
    if (io_en) begin
      o3 <= o2;
    end
    if (io_en) begin
      o4 <= o3;
    end
    if (io_en) begin
      r5 <= _T_4;
    end
    if (io_en) begin
      r6 <= r5;
    end
  end
endmodule
module Loaf(
  input         clock,
  input         reset,
  input         io_start,
  output        io_doneLoading,
  input         io_modeLoad,
  input         io_modeCompute,
  input         io_loadIdx,
  input         io_computeIdx,
  output        io_off_ready,
  input         io_off_valid,
  input  [15:0] io_off_bits_0,
  input  [15:0] io_off_bits_1,
  input  [15:0] io_off_bits_2,
  input  [15:0] io_off_bits_3,
  input  [15:0] io_off_bits_4,
  input  [15:0] io_off_bits_5,
  input  [15:0] io_off_bits_6,
  input  [15:0] io_off_bits_7,
  input         io_out_ready,
  output        io_out_valid,
  output [15:0] io_out_bits_0,
  output [15:0] io_out_bits_1,
  output [15:0] io_out_bits_2,
  output [15:0] io_out_bits_3,
  output [15:0] io_out_bits_4,
  output [15:0] io_out_bits_5,
  output [15:0] io_out_bits_6,
  output [15:0] io_out_bits_7,
  output        io_slc_ready,
  input         io_slc_valid,
  input  [15:0] io_slc_bits_e,
  input  [15:0] io_slc_bits_a,
  output        io_lof_ready,
  input         io_lof_valid,
  input  [15:0] io_lof_bits_e,
  input  [15:0] io_lof_bits_a
);
  wire  macs_0_0_clock; // @[loaf.scala 120:72]
  wire  macs_0_0_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_0_0_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_0_0_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_0_0_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_0_0_io_r; // @[loaf.scala 120:72]
  wire  macs_0_1_clock; // @[loaf.scala 120:72]
  wire  macs_0_1_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_0_1_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_0_1_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_0_1_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_0_1_io_r; // @[loaf.scala 120:72]
  wire  macs_0_2_clock; // @[loaf.scala 120:72]
  wire  macs_0_2_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_0_2_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_0_2_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_0_2_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_0_2_io_r; // @[loaf.scala 120:72]
  wire  macs_0_3_clock; // @[loaf.scala 120:72]
  wire  macs_0_3_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_0_3_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_0_3_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_0_3_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_0_3_io_r; // @[loaf.scala 120:72]
  wire  macs_0_4_clock; // @[loaf.scala 120:72]
  wire  macs_0_4_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_0_4_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_0_4_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_0_4_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_0_4_io_r; // @[loaf.scala 120:72]
  wire  macs_0_5_clock; // @[loaf.scala 120:72]
  wire  macs_0_5_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_0_5_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_0_5_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_0_5_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_0_5_io_r; // @[loaf.scala 120:72]
  wire  macs_0_6_clock; // @[loaf.scala 120:72]
  wire  macs_0_6_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_0_6_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_0_6_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_0_6_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_0_6_io_r; // @[loaf.scala 120:72]
  wire  macs_0_7_clock; // @[loaf.scala 120:72]
  wire  macs_0_7_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_0_7_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_0_7_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_0_7_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_0_7_io_r; // @[loaf.scala 120:72]
  wire  macs_1_0_clock; // @[loaf.scala 120:72]
  wire  macs_1_0_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_1_0_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_1_0_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_1_0_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_1_0_io_r; // @[loaf.scala 120:72]
  wire  macs_1_1_clock; // @[loaf.scala 120:72]
  wire  macs_1_1_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_1_1_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_1_1_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_1_1_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_1_1_io_r; // @[loaf.scala 120:72]
  wire  macs_1_2_clock; // @[loaf.scala 120:72]
  wire  macs_1_2_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_1_2_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_1_2_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_1_2_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_1_2_io_r; // @[loaf.scala 120:72]
  wire  macs_1_3_clock; // @[loaf.scala 120:72]
  wire  macs_1_3_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_1_3_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_1_3_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_1_3_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_1_3_io_r; // @[loaf.scala 120:72]
  wire  macs_1_4_clock; // @[loaf.scala 120:72]
  wire  macs_1_4_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_1_4_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_1_4_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_1_4_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_1_4_io_r; // @[loaf.scala 120:72]
  wire  macs_1_5_clock; // @[loaf.scala 120:72]
  wire  macs_1_5_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_1_5_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_1_5_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_1_5_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_1_5_io_r; // @[loaf.scala 120:72]
  wire  macs_1_6_clock; // @[loaf.scala 120:72]
  wire  macs_1_6_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_1_6_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_1_6_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_1_6_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_1_6_io_r; // @[loaf.scala 120:72]
  wire  macs_1_7_clock; // @[loaf.scala 120:72]
  wire  macs_1_7_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_1_7_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_1_7_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_1_7_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_1_7_io_r; // @[loaf.scala 120:72]
  wire  macs_2_0_clock; // @[loaf.scala 120:72]
  wire  macs_2_0_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_2_0_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_2_0_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_2_0_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_2_0_io_r; // @[loaf.scala 120:72]
  wire  macs_2_1_clock; // @[loaf.scala 120:72]
  wire  macs_2_1_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_2_1_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_2_1_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_2_1_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_2_1_io_r; // @[loaf.scala 120:72]
  wire  macs_2_2_clock; // @[loaf.scala 120:72]
  wire  macs_2_2_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_2_2_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_2_2_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_2_2_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_2_2_io_r; // @[loaf.scala 120:72]
  wire  macs_2_3_clock; // @[loaf.scala 120:72]
  wire  macs_2_3_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_2_3_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_2_3_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_2_3_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_2_3_io_r; // @[loaf.scala 120:72]
  wire  macs_2_4_clock; // @[loaf.scala 120:72]
  wire  macs_2_4_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_2_4_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_2_4_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_2_4_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_2_4_io_r; // @[loaf.scala 120:72]
  wire  macs_2_5_clock; // @[loaf.scala 120:72]
  wire  macs_2_5_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_2_5_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_2_5_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_2_5_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_2_5_io_r; // @[loaf.scala 120:72]
  wire  macs_2_6_clock; // @[loaf.scala 120:72]
  wire  macs_2_6_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_2_6_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_2_6_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_2_6_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_2_6_io_r; // @[loaf.scala 120:72]
  wire  macs_2_7_clock; // @[loaf.scala 120:72]
  wire  macs_2_7_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_2_7_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_2_7_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_2_7_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_2_7_io_r; // @[loaf.scala 120:72]
  wire  macs_3_0_clock; // @[loaf.scala 120:72]
  wire  macs_3_0_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_3_0_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_3_0_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_3_0_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_3_0_io_r; // @[loaf.scala 120:72]
  wire  macs_3_1_clock; // @[loaf.scala 120:72]
  wire  macs_3_1_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_3_1_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_3_1_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_3_1_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_3_1_io_r; // @[loaf.scala 120:72]
  wire  macs_3_2_clock; // @[loaf.scala 120:72]
  wire  macs_3_2_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_3_2_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_3_2_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_3_2_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_3_2_io_r; // @[loaf.scala 120:72]
  wire  macs_3_3_clock; // @[loaf.scala 120:72]
  wire  macs_3_3_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_3_3_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_3_3_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_3_3_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_3_3_io_r; // @[loaf.scala 120:72]
  wire  macs_3_4_clock; // @[loaf.scala 120:72]
  wire  macs_3_4_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_3_4_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_3_4_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_3_4_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_3_4_io_r; // @[loaf.scala 120:72]
  wire  macs_3_5_clock; // @[loaf.scala 120:72]
  wire  macs_3_5_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_3_5_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_3_5_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_3_5_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_3_5_io_r; // @[loaf.scala 120:72]
  wire  macs_3_6_clock; // @[loaf.scala 120:72]
  wire  macs_3_6_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_3_6_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_3_6_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_3_6_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_3_6_io_r; // @[loaf.scala 120:72]
  wire  macs_3_7_clock; // @[loaf.scala 120:72]
  wire  macs_3_7_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_3_7_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_3_7_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_3_7_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_3_7_io_r; // @[loaf.scala 120:72]
  wire  macs_4_0_clock; // @[loaf.scala 120:72]
  wire  macs_4_0_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_4_0_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_4_0_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_4_0_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_4_0_io_r; // @[loaf.scala 120:72]
  wire  macs_4_1_clock; // @[loaf.scala 120:72]
  wire  macs_4_1_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_4_1_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_4_1_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_4_1_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_4_1_io_r; // @[loaf.scala 120:72]
  wire  macs_4_2_clock; // @[loaf.scala 120:72]
  wire  macs_4_2_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_4_2_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_4_2_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_4_2_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_4_2_io_r; // @[loaf.scala 120:72]
  wire  macs_4_3_clock; // @[loaf.scala 120:72]
  wire  macs_4_3_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_4_3_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_4_3_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_4_3_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_4_3_io_r; // @[loaf.scala 120:72]
  wire  macs_4_4_clock; // @[loaf.scala 120:72]
  wire  macs_4_4_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_4_4_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_4_4_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_4_4_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_4_4_io_r; // @[loaf.scala 120:72]
  wire  macs_4_5_clock; // @[loaf.scala 120:72]
  wire  macs_4_5_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_4_5_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_4_5_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_4_5_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_4_5_io_r; // @[loaf.scala 120:72]
  wire  macs_4_6_clock; // @[loaf.scala 120:72]
  wire  macs_4_6_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_4_6_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_4_6_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_4_6_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_4_6_io_r; // @[loaf.scala 120:72]
  wire  macs_4_7_clock; // @[loaf.scala 120:72]
  wire  macs_4_7_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_4_7_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_4_7_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_4_7_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_4_7_io_r; // @[loaf.scala 120:72]
  wire  macs_5_0_clock; // @[loaf.scala 120:72]
  wire  macs_5_0_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_5_0_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_5_0_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_5_0_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_5_0_io_r; // @[loaf.scala 120:72]
  wire  macs_5_1_clock; // @[loaf.scala 120:72]
  wire  macs_5_1_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_5_1_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_5_1_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_5_1_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_5_1_io_r; // @[loaf.scala 120:72]
  wire  macs_5_2_clock; // @[loaf.scala 120:72]
  wire  macs_5_2_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_5_2_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_5_2_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_5_2_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_5_2_io_r; // @[loaf.scala 120:72]
  wire  macs_5_3_clock; // @[loaf.scala 120:72]
  wire  macs_5_3_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_5_3_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_5_3_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_5_3_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_5_3_io_r; // @[loaf.scala 120:72]
  wire  macs_5_4_clock; // @[loaf.scala 120:72]
  wire  macs_5_4_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_5_4_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_5_4_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_5_4_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_5_4_io_r; // @[loaf.scala 120:72]
  wire  macs_5_5_clock; // @[loaf.scala 120:72]
  wire  macs_5_5_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_5_5_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_5_5_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_5_5_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_5_5_io_r; // @[loaf.scala 120:72]
  wire  macs_5_6_clock; // @[loaf.scala 120:72]
  wire  macs_5_6_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_5_6_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_5_6_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_5_6_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_5_6_io_r; // @[loaf.scala 120:72]
  wire  macs_5_7_clock; // @[loaf.scala 120:72]
  wire  macs_5_7_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_5_7_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_5_7_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_5_7_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_5_7_io_r; // @[loaf.scala 120:72]
  wire  macs_6_0_clock; // @[loaf.scala 120:72]
  wire  macs_6_0_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_6_0_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_6_0_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_6_0_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_6_0_io_r; // @[loaf.scala 120:72]
  wire  macs_6_1_clock; // @[loaf.scala 120:72]
  wire  macs_6_1_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_6_1_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_6_1_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_6_1_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_6_1_io_r; // @[loaf.scala 120:72]
  wire  macs_6_2_clock; // @[loaf.scala 120:72]
  wire  macs_6_2_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_6_2_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_6_2_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_6_2_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_6_2_io_r; // @[loaf.scala 120:72]
  wire  macs_6_3_clock; // @[loaf.scala 120:72]
  wire  macs_6_3_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_6_3_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_6_3_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_6_3_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_6_3_io_r; // @[loaf.scala 120:72]
  wire  macs_6_4_clock; // @[loaf.scala 120:72]
  wire  macs_6_4_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_6_4_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_6_4_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_6_4_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_6_4_io_r; // @[loaf.scala 120:72]
  wire  macs_6_5_clock; // @[loaf.scala 120:72]
  wire  macs_6_5_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_6_5_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_6_5_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_6_5_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_6_5_io_r; // @[loaf.scala 120:72]
  wire  macs_6_6_clock; // @[loaf.scala 120:72]
  wire  macs_6_6_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_6_6_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_6_6_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_6_6_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_6_6_io_r; // @[loaf.scala 120:72]
  wire  macs_6_7_clock; // @[loaf.scala 120:72]
  wire  macs_6_7_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_6_7_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_6_7_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_6_7_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_6_7_io_r; // @[loaf.scala 120:72]
  wire  macs_7_0_clock; // @[loaf.scala 120:72]
  wire  macs_7_0_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_7_0_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_7_0_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_7_0_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_7_0_io_r; // @[loaf.scala 120:72]
  wire  macs_7_1_clock; // @[loaf.scala 120:72]
  wire  macs_7_1_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_7_1_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_7_1_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_7_1_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_7_1_io_r; // @[loaf.scala 120:72]
  wire  macs_7_2_clock; // @[loaf.scala 120:72]
  wire  macs_7_2_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_7_2_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_7_2_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_7_2_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_7_2_io_r; // @[loaf.scala 120:72]
  wire  macs_7_3_clock; // @[loaf.scala 120:72]
  wire  macs_7_3_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_7_3_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_7_3_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_7_3_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_7_3_io_r; // @[loaf.scala 120:72]
  wire  macs_7_4_clock; // @[loaf.scala 120:72]
  wire  macs_7_4_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_7_4_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_7_4_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_7_4_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_7_4_io_r; // @[loaf.scala 120:72]
  wire  macs_7_5_clock; // @[loaf.scala 120:72]
  wire  macs_7_5_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_7_5_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_7_5_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_7_5_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_7_5_io_r; // @[loaf.scala 120:72]
  wire  macs_7_6_clock; // @[loaf.scala 120:72]
  wire  macs_7_6_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_7_6_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_7_6_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_7_6_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_7_6_io_r; // @[loaf.scala 120:72]
  wire  macs_7_7_clock; // @[loaf.scala 120:72]
  wire  macs_7_7_io_en; // @[loaf.scala 120:72]
  wire [15:0] macs_7_7_io_a; // @[loaf.scala 120:72]
  wire [15:0] macs_7_7_io_b; // @[loaf.scala 120:72]
  wire [31:0] macs_7_7_io_o; // @[loaf.scala 120:72]
  wire [31:0] macs_7_7_io_r; // @[loaf.scala 120:72]
  reg [31:0] AE_0_0 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_0;
  wire [31:0] AE_0_0__T_497_data; // @[loaf.scala 147:67]
  wire [4:0] AE_0_0__T_497_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_0_0__T_9_data; // @[loaf.scala 147:67]
  wire [4:0] AE_0_0__T_9_addr; // @[loaf.scala 147:67]
  wire  AE_0_0__T_9_mask; // @[loaf.scala 147:67]
  wire  AE_0_0__T_9_en; // @[loaf.scala 147:67]
  reg [31:0] AE_0_1 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_1;
  wire [31:0] AE_0_1__T_585_data; // @[loaf.scala 147:67]
  wire [4:0] AE_0_1__T_585_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_0_1__T_15_data; // @[loaf.scala 147:67]
  wire [4:0] AE_0_1__T_15_addr; // @[loaf.scala 147:67]
  wire  AE_0_1__T_15_mask; // @[loaf.scala 147:67]
  wire  AE_0_1__T_15_en; // @[loaf.scala 147:67]
  reg [31:0] AE_0_2 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_2;
  wire [31:0] AE_0_2__T_673_data; // @[loaf.scala 147:67]
  wire [4:0] AE_0_2__T_673_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_0_2__T_21_data; // @[loaf.scala 147:67]
  wire [4:0] AE_0_2__T_21_addr; // @[loaf.scala 147:67]
  wire  AE_0_2__T_21_mask; // @[loaf.scala 147:67]
  wire  AE_0_2__T_21_en; // @[loaf.scala 147:67]
  reg [31:0] AE_0_3 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_3;
  wire [31:0] AE_0_3__T_761_data; // @[loaf.scala 147:67]
  wire [4:0] AE_0_3__T_761_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_0_3__T_27_data; // @[loaf.scala 147:67]
  wire [4:0] AE_0_3__T_27_addr; // @[loaf.scala 147:67]
  wire  AE_0_3__T_27_mask; // @[loaf.scala 147:67]
  wire  AE_0_3__T_27_en; // @[loaf.scala 147:67]
  reg [31:0] AE_0_4 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_4;
  wire [31:0] AE_0_4__T_849_data; // @[loaf.scala 147:67]
  wire [4:0] AE_0_4__T_849_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_0_4__T_33_data; // @[loaf.scala 147:67]
  wire [4:0] AE_0_4__T_33_addr; // @[loaf.scala 147:67]
  wire  AE_0_4__T_33_mask; // @[loaf.scala 147:67]
  wire  AE_0_4__T_33_en; // @[loaf.scala 147:67]
  reg [31:0] AE_0_5 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_5;
  wire [31:0] AE_0_5__T_937_data; // @[loaf.scala 147:67]
  wire [4:0] AE_0_5__T_937_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_0_5__T_39_data; // @[loaf.scala 147:67]
  wire [4:0] AE_0_5__T_39_addr; // @[loaf.scala 147:67]
  wire  AE_0_5__T_39_mask; // @[loaf.scala 147:67]
  wire  AE_0_5__T_39_en; // @[loaf.scala 147:67]
  reg [31:0] AE_0_6 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_6;
  wire [31:0] AE_0_6__T_1025_data; // @[loaf.scala 147:67]
  wire [4:0] AE_0_6__T_1025_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_0_6__T_45_data; // @[loaf.scala 147:67]
  wire [4:0] AE_0_6__T_45_addr; // @[loaf.scala 147:67]
  wire  AE_0_6__T_45_mask; // @[loaf.scala 147:67]
  wire  AE_0_6__T_45_en; // @[loaf.scala 147:67]
  reg [31:0] AE_0_7 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_7;
  wire [31:0] AE_0_7__T_1113_data; // @[loaf.scala 147:67]
  wire [4:0] AE_0_7__T_1113_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_0_7__T_51_data; // @[loaf.scala 147:67]
  wire [4:0] AE_0_7__T_51_addr; // @[loaf.scala 147:67]
  wire  AE_0_7__T_51_mask; // @[loaf.scala 147:67]
  wire  AE_0_7__T_51_en; // @[loaf.scala 147:67]
  reg [31:0] AE_1_0 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_8;
  wire [31:0] AE_1_0__T_508_data; // @[loaf.scala 147:67]
  wire [4:0] AE_1_0__T_508_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_1_0__T_57_data; // @[loaf.scala 147:67]
  wire [4:0] AE_1_0__T_57_addr; // @[loaf.scala 147:67]
  wire  AE_1_0__T_57_mask; // @[loaf.scala 147:67]
  wire  AE_1_0__T_57_en; // @[loaf.scala 147:67]
  reg [31:0] AE_1_1 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_9;
  wire [31:0] AE_1_1__T_596_data; // @[loaf.scala 147:67]
  wire [4:0] AE_1_1__T_596_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_1_1__T_63_data; // @[loaf.scala 147:67]
  wire [4:0] AE_1_1__T_63_addr; // @[loaf.scala 147:67]
  wire  AE_1_1__T_63_mask; // @[loaf.scala 147:67]
  wire  AE_1_1__T_63_en; // @[loaf.scala 147:67]
  reg [31:0] AE_1_2 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_10;
  wire [31:0] AE_1_2__T_684_data; // @[loaf.scala 147:67]
  wire [4:0] AE_1_2__T_684_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_1_2__T_69_data; // @[loaf.scala 147:67]
  wire [4:0] AE_1_2__T_69_addr; // @[loaf.scala 147:67]
  wire  AE_1_2__T_69_mask; // @[loaf.scala 147:67]
  wire  AE_1_2__T_69_en; // @[loaf.scala 147:67]
  reg [31:0] AE_1_3 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_11;
  wire [31:0] AE_1_3__T_772_data; // @[loaf.scala 147:67]
  wire [4:0] AE_1_3__T_772_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_1_3__T_75_data; // @[loaf.scala 147:67]
  wire [4:0] AE_1_3__T_75_addr; // @[loaf.scala 147:67]
  wire  AE_1_3__T_75_mask; // @[loaf.scala 147:67]
  wire  AE_1_3__T_75_en; // @[loaf.scala 147:67]
  reg [31:0] AE_1_4 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_12;
  wire [31:0] AE_1_4__T_860_data; // @[loaf.scala 147:67]
  wire [4:0] AE_1_4__T_860_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_1_4__T_81_data; // @[loaf.scala 147:67]
  wire [4:0] AE_1_4__T_81_addr; // @[loaf.scala 147:67]
  wire  AE_1_4__T_81_mask; // @[loaf.scala 147:67]
  wire  AE_1_4__T_81_en; // @[loaf.scala 147:67]
  reg [31:0] AE_1_5 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_13;
  wire [31:0] AE_1_5__T_948_data; // @[loaf.scala 147:67]
  wire [4:0] AE_1_5__T_948_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_1_5__T_87_data; // @[loaf.scala 147:67]
  wire [4:0] AE_1_5__T_87_addr; // @[loaf.scala 147:67]
  wire  AE_1_5__T_87_mask; // @[loaf.scala 147:67]
  wire  AE_1_5__T_87_en; // @[loaf.scala 147:67]
  reg [31:0] AE_1_6 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_14;
  wire [31:0] AE_1_6__T_1036_data; // @[loaf.scala 147:67]
  wire [4:0] AE_1_6__T_1036_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_1_6__T_93_data; // @[loaf.scala 147:67]
  wire [4:0] AE_1_6__T_93_addr; // @[loaf.scala 147:67]
  wire  AE_1_6__T_93_mask; // @[loaf.scala 147:67]
  wire  AE_1_6__T_93_en; // @[loaf.scala 147:67]
  reg [31:0] AE_1_7 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_15;
  wire [31:0] AE_1_7__T_1124_data; // @[loaf.scala 147:67]
  wire [4:0] AE_1_7__T_1124_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_1_7__T_99_data; // @[loaf.scala 147:67]
  wire [4:0] AE_1_7__T_99_addr; // @[loaf.scala 147:67]
  wire  AE_1_7__T_99_mask; // @[loaf.scala 147:67]
  wire  AE_1_7__T_99_en; // @[loaf.scala 147:67]
  reg [31:0] AE_2_0 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_16;
  wire [31:0] AE_2_0__T_519_data; // @[loaf.scala 147:67]
  wire [4:0] AE_2_0__T_519_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_2_0__T_105_data; // @[loaf.scala 147:67]
  wire [4:0] AE_2_0__T_105_addr; // @[loaf.scala 147:67]
  wire  AE_2_0__T_105_mask; // @[loaf.scala 147:67]
  wire  AE_2_0__T_105_en; // @[loaf.scala 147:67]
  reg [31:0] AE_2_1 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_17;
  wire [31:0] AE_2_1__T_607_data; // @[loaf.scala 147:67]
  wire [4:0] AE_2_1__T_607_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_2_1__T_111_data; // @[loaf.scala 147:67]
  wire [4:0] AE_2_1__T_111_addr; // @[loaf.scala 147:67]
  wire  AE_2_1__T_111_mask; // @[loaf.scala 147:67]
  wire  AE_2_1__T_111_en; // @[loaf.scala 147:67]
  reg [31:0] AE_2_2 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_18;
  wire [31:0] AE_2_2__T_695_data; // @[loaf.scala 147:67]
  wire [4:0] AE_2_2__T_695_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_2_2__T_117_data; // @[loaf.scala 147:67]
  wire [4:0] AE_2_2__T_117_addr; // @[loaf.scala 147:67]
  wire  AE_2_2__T_117_mask; // @[loaf.scala 147:67]
  wire  AE_2_2__T_117_en; // @[loaf.scala 147:67]
  reg [31:0] AE_2_3 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_19;
  wire [31:0] AE_2_3__T_783_data; // @[loaf.scala 147:67]
  wire [4:0] AE_2_3__T_783_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_2_3__T_123_data; // @[loaf.scala 147:67]
  wire [4:0] AE_2_3__T_123_addr; // @[loaf.scala 147:67]
  wire  AE_2_3__T_123_mask; // @[loaf.scala 147:67]
  wire  AE_2_3__T_123_en; // @[loaf.scala 147:67]
  reg [31:0] AE_2_4 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_20;
  wire [31:0] AE_2_4__T_871_data; // @[loaf.scala 147:67]
  wire [4:0] AE_2_4__T_871_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_2_4__T_129_data; // @[loaf.scala 147:67]
  wire [4:0] AE_2_4__T_129_addr; // @[loaf.scala 147:67]
  wire  AE_2_4__T_129_mask; // @[loaf.scala 147:67]
  wire  AE_2_4__T_129_en; // @[loaf.scala 147:67]
  reg [31:0] AE_2_5 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_21;
  wire [31:0] AE_2_5__T_959_data; // @[loaf.scala 147:67]
  wire [4:0] AE_2_5__T_959_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_2_5__T_135_data; // @[loaf.scala 147:67]
  wire [4:0] AE_2_5__T_135_addr; // @[loaf.scala 147:67]
  wire  AE_2_5__T_135_mask; // @[loaf.scala 147:67]
  wire  AE_2_5__T_135_en; // @[loaf.scala 147:67]
  reg [31:0] AE_2_6 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_22;
  wire [31:0] AE_2_6__T_1047_data; // @[loaf.scala 147:67]
  wire [4:0] AE_2_6__T_1047_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_2_6__T_141_data; // @[loaf.scala 147:67]
  wire [4:0] AE_2_6__T_141_addr; // @[loaf.scala 147:67]
  wire  AE_2_6__T_141_mask; // @[loaf.scala 147:67]
  wire  AE_2_6__T_141_en; // @[loaf.scala 147:67]
  reg [31:0] AE_2_7 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_23;
  wire [31:0] AE_2_7__T_1135_data; // @[loaf.scala 147:67]
  wire [4:0] AE_2_7__T_1135_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_2_7__T_147_data; // @[loaf.scala 147:67]
  wire [4:0] AE_2_7__T_147_addr; // @[loaf.scala 147:67]
  wire  AE_2_7__T_147_mask; // @[loaf.scala 147:67]
  wire  AE_2_7__T_147_en; // @[loaf.scala 147:67]
  reg [31:0] AE_3_0 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_24;
  wire [31:0] AE_3_0__T_530_data; // @[loaf.scala 147:67]
  wire [4:0] AE_3_0__T_530_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_3_0__T_153_data; // @[loaf.scala 147:67]
  wire [4:0] AE_3_0__T_153_addr; // @[loaf.scala 147:67]
  wire  AE_3_0__T_153_mask; // @[loaf.scala 147:67]
  wire  AE_3_0__T_153_en; // @[loaf.scala 147:67]
  reg [31:0] AE_3_1 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_25;
  wire [31:0] AE_3_1__T_618_data; // @[loaf.scala 147:67]
  wire [4:0] AE_3_1__T_618_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_3_1__T_159_data; // @[loaf.scala 147:67]
  wire [4:0] AE_3_1__T_159_addr; // @[loaf.scala 147:67]
  wire  AE_3_1__T_159_mask; // @[loaf.scala 147:67]
  wire  AE_3_1__T_159_en; // @[loaf.scala 147:67]
  reg [31:0] AE_3_2 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_26;
  wire [31:0] AE_3_2__T_706_data; // @[loaf.scala 147:67]
  wire [4:0] AE_3_2__T_706_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_3_2__T_165_data; // @[loaf.scala 147:67]
  wire [4:0] AE_3_2__T_165_addr; // @[loaf.scala 147:67]
  wire  AE_3_2__T_165_mask; // @[loaf.scala 147:67]
  wire  AE_3_2__T_165_en; // @[loaf.scala 147:67]
  reg [31:0] AE_3_3 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_27;
  wire [31:0] AE_3_3__T_794_data; // @[loaf.scala 147:67]
  wire [4:0] AE_3_3__T_794_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_3_3__T_171_data; // @[loaf.scala 147:67]
  wire [4:0] AE_3_3__T_171_addr; // @[loaf.scala 147:67]
  wire  AE_3_3__T_171_mask; // @[loaf.scala 147:67]
  wire  AE_3_3__T_171_en; // @[loaf.scala 147:67]
  reg [31:0] AE_3_4 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_28;
  wire [31:0] AE_3_4__T_882_data; // @[loaf.scala 147:67]
  wire [4:0] AE_3_4__T_882_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_3_4__T_177_data; // @[loaf.scala 147:67]
  wire [4:0] AE_3_4__T_177_addr; // @[loaf.scala 147:67]
  wire  AE_3_4__T_177_mask; // @[loaf.scala 147:67]
  wire  AE_3_4__T_177_en; // @[loaf.scala 147:67]
  reg [31:0] AE_3_5 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_29;
  wire [31:0] AE_3_5__T_970_data; // @[loaf.scala 147:67]
  wire [4:0] AE_3_5__T_970_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_3_5__T_183_data; // @[loaf.scala 147:67]
  wire [4:0] AE_3_5__T_183_addr; // @[loaf.scala 147:67]
  wire  AE_3_5__T_183_mask; // @[loaf.scala 147:67]
  wire  AE_3_5__T_183_en; // @[loaf.scala 147:67]
  reg [31:0] AE_3_6 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_30;
  wire [31:0] AE_3_6__T_1058_data; // @[loaf.scala 147:67]
  wire [4:0] AE_3_6__T_1058_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_3_6__T_189_data; // @[loaf.scala 147:67]
  wire [4:0] AE_3_6__T_189_addr; // @[loaf.scala 147:67]
  wire  AE_3_6__T_189_mask; // @[loaf.scala 147:67]
  wire  AE_3_6__T_189_en; // @[loaf.scala 147:67]
  reg [31:0] AE_3_7 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_31;
  wire [31:0] AE_3_7__T_1146_data; // @[loaf.scala 147:67]
  wire [4:0] AE_3_7__T_1146_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_3_7__T_195_data; // @[loaf.scala 147:67]
  wire [4:0] AE_3_7__T_195_addr; // @[loaf.scala 147:67]
  wire  AE_3_7__T_195_mask; // @[loaf.scala 147:67]
  wire  AE_3_7__T_195_en; // @[loaf.scala 147:67]
  reg [31:0] AE_4_0 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_32;
  wire [31:0] AE_4_0__T_541_data; // @[loaf.scala 147:67]
  wire [4:0] AE_4_0__T_541_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_4_0__T_201_data; // @[loaf.scala 147:67]
  wire [4:0] AE_4_0__T_201_addr; // @[loaf.scala 147:67]
  wire  AE_4_0__T_201_mask; // @[loaf.scala 147:67]
  wire  AE_4_0__T_201_en; // @[loaf.scala 147:67]
  reg [31:0] AE_4_1 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_33;
  wire [31:0] AE_4_1__T_629_data; // @[loaf.scala 147:67]
  wire [4:0] AE_4_1__T_629_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_4_1__T_207_data; // @[loaf.scala 147:67]
  wire [4:0] AE_4_1__T_207_addr; // @[loaf.scala 147:67]
  wire  AE_4_1__T_207_mask; // @[loaf.scala 147:67]
  wire  AE_4_1__T_207_en; // @[loaf.scala 147:67]
  reg [31:0] AE_4_2 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_34;
  wire [31:0] AE_4_2__T_717_data; // @[loaf.scala 147:67]
  wire [4:0] AE_4_2__T_717_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_4_2__T_213_data; // @[loaf.scala 147:67]
  wire [4:0] AE_4_2__T_213_addr; // @[loaf.scala 147:67]
  wire  AE_4_2__T_213_mask; // @[loaf.scala 147:67]
  wire  AE_4_2__T_213_en; // @[loaf.scala 147:67]
  reg [31:0] AE_4_3 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_35;
  wire [31:0] AE_4_3__T_805_data; // @[loaf.scala 147:67]
  wire [4:0] AE_4_3__T_805_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_4_3__T_219_data; // @[loaf.scala 147:67]
  wire [4:0] AE_4_3__T_219_addr; // @[loaf.scala 147:67]
  wire  AE_4_3__T_219_mask; // @[loaf.scala 147:67]
  wire  AE_4_3__T_219_en; // @[loaf.scala 147:67]
  reg [31:0] AE_4_4 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_36;
  wire [31:0] AE_4_4__T_893_data; // @[loaf.scala 147:67]
  wire [4:0] AE_4_4__T_893_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_4_4__T_225_data; // @[loaf.scala 147:67]
  wire [4:0] AE_4_4__T_225_addr; // @[loaf.scala 147:67]
  wire  AE_4_4__T_225_mask; // @[loaf.scala 147:67]
  wire  AE_4_4__T_225_en; // @[loaf.scala 147:67]
  reg [31:0] AE_4_5 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_37;
  wire [31:0] AE_4_5__T_981_data; // @[loaf.scala 147:67]
  wire [4:0] AE_4_5__T_981_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_4_5__T_231_data; // @[loaf.scala 147:67]
  wire [4:0] AE_4_5__T_231_addr; // @[loaf.scala 147:67]
  wire  AE_4_5__T_231_mask; // @[loaf.scala 147:67]
  wire  AE_4_5__T_231_en; // @[loaf.scala 147:67]
  reg [31:0] AE_4_6 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_38;
  wire [31:0] AE_4_6__T_1069_data; // @[loaf.scala 147:67]
  wire [4:0] AE_4_6__T_1069_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_4_6__T_237_data; // @[loaf.scala 147:67]
  wire [4:0] AE_4_6__T_237_addr; // @[loaf.scala 147:67]
  wire  AE_4_6__T_237_mask; // @[loaf.scala 147:67]
  wire  AE_4_6__T_237_en; // @[loaf.scala 147:67]
  reg [31:0] AE_4_7 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_39;
  wire [31:0] AE_4_7__T_1157_data; // @[loaf.scala 147:67]
  wire [4:0] AE_4_7__T_1157_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_4_7__T_243_data; // @[loaf.scala 147:67]
  wire [4:0] AE_4_7__T_243_addr; // @[loaf.scala 147:67]
  wire  AE_4_7__T_243_mask; // @[loaf.scala 147:67]
  wire  AE_4_7__T_243_en; // @[loaf.scala 147:67]
  reg [31:0] AE_5_0 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_40;
  wire [31:0] AE_5_0__T_552_data; // @[loaf.scala 147:67]
  wire [4:0] AE_5_0__T_552_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_5_0__T_249_data; // @[loaf.scala 147:67]
  wire [4:0] AE_5_0__T_249_addr; // @[loaf.scala 147:67]
  wire  AE_5_0__T_249_mask; // @[loaf.scala 147:67]
  wire  AE_5_0__T_249_en; // @[loaf.scala 147:67]
  reg [31:0] AE_5_1 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_41;
  wire [31:0] AE_5_1__T_640_data; // @[loaf.scala 147:67]
  wire [4:0] AE_5_1__T_640_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_5_1__T_255_data; // @[loaf.scala 147:67]
  wire [4:0] AE_5_1__T_255_addr; // @[loaf.scala 147:67]
  wire  AE_5_1__T_255_mask; // @[loaf.scala 147:67]
  wire  AE_5_1__T_255_en; // @[loaf.scala 147:67]
  reg [31:0] AE_5_2 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_42;
  wire [31:0] AE_5_2__T_728_data; // @[loaf.scala 147:67]
  wire [4:0] AE_5_2__T_728_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_5_2__T_261_data; // @[loaf.scala 147:67]
  wire [4:0] AE_5_2__T_261_addr; // @[loaf.scala 147:67]
  wire  AE_5_2__T_261_mask; // @[loaf.scala 147:67]
  wire  AE_5_2__T_261_en; // @[loaf.scala 147:67]
  reg [31:0] AE_5_3 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_43;
  wire [31:0] AE_5_3__T_816_data; // @[loaf.scala 147:67]
  wire [4:0] AE_5_3__T_816_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_5_3__T_267_data; // @[loaf.scala 147:67]
  wire [4:0] AE_5_3__T_267_addr; // @[loaf.scala 147:67]
  wire  AE_5_3__T_267_mask; // @[loaf.scala 147:67]
  wire  AE_5_3__T_267_en; // @[loaf.scala 147:67]
  reg [31:0] AE_5_4 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_44;
  wire [31:0] AE_5_4__T_904_data; // @[loaf.scala 147:67]
  wire [4:0] AE_5_4__T_904_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_5_4__T_273_data; // @[loaf.scala 147:67]
  wire [4:0] AE_5_4__T_273_addr; // @[loaf.scala 147:67]
  wire  AE_5_4__T_273_mask; // @[loaf.scala 147:67]
  wire  AE_5_4__T_273_en; // @[loaf.scala 147:67]
  reg [31:0] AE_5_5 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_45;
  wire [31:0] AE_5_5__T_992_data; // @[loaf.scala 147:67]
  wire [4:0] AE_5_5__T_992_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_5_5__T_279_data; // @[loaf.scala 147:67]
  wire [4:0] AE_5_5__T_279_addr; // @[loaf.scala 147:67]
  wire  AE_5_5__T_279_mask; // @[loaf.scala 147:67]
  wire  AE_5_5__T_279_en; // @[loaf.scala 147:67]
  reg [31:0] AE_5_6 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_46;
  wire [31:0] AE_5_6__T_1080_data; // @[loaf.scala 147:67]
  wire [4:0] AE_5_6__T_1080_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_5_6__T_285_data; // @[loaf.scala 147:67]
  wire [4:0] AE_5_6__T_285_addr; // @[loaf.scala 147:67]
  wire  AE_5_6__T_285_mask; // @[loaf.scala 147:67]
  wire  AE_5_6__T_285_en; // @[loaf.scala 147:67]
  reg [31:0] AE_5_7 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_47;
  wire [31:0] AE_5_7__T_1168_data; // @[loaf.scala 147:67]
  wire [4:0] AE_5_7__T_1168_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_5_7__T_291_data; // @[loaf.scala 147:67]
  wire [4:0] AE_5_7__T_291_addr; // @[loaf.scala 147:67]
  wire  AE_5_7__T_291_mask; // @[loaf.scala 147:67]
  wire  AE_5_7__T_291_en; // @[loaf.scala 147:67]
  reg [31:0] AE_6_0 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_48;
  wire [31:0] AE_6_0__T_563_data; // @[loaf.scala 147:67]
  wire [4:0] AE_6_0__T_563_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_6_0__T_297_data; // @[loaf.scala 147:67]
  wire [4:0] AE_6_0__T_297_addr; // @[loaf.scala 147:67]
  wire  AE_6_0__T_297_mask; // @[loaf.scala 147:67]
  wire  AE_6_0__T_297_en; // @[loaf.scala 147:67]
  reg [31:0] AE_6_1 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_49;
  wire [31:0] AE_6_1__T_651_data; // @[loaf.scala 147:67]
  wire [4:0] AE_6_1__T_651_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_6_1__T_303_data; // @[loaf.scala 147:67]
  wire [4:0] AE_6_1__T_303_addr; // @[loaf.scala 147:67]
  wire  AE_6_1__T_303_mask; // @[loaf.scala 147:67]
  wire  AE_6_1__T_303_en; // @[loaf.scala 147:67]
  reg [31:0] AE_6_2 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_50;
  wire [31:0] AE_6_2__T_739_data; // @[loaf.scala 147:67]
  wire [4:0] AE_6_2__T_739_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_6_2__T_309_data; // @[loaf.scala 147:67]
  wire [4:0] AE_6_2__T_309_addr; // @[loaf.scala 147:67]
  wire  AE_6_2__T_309_mask; // @[loaf.scala 147:67]
  wire  AE_6_2__T_309_en; // @[loaf.scala 147:67]
  reg [31:0] AE_6_3 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_51;
  wire [31:0] AE_6_3__T_827_data; // @[loaf.scala 147:67]
  wire [4:0] AE_6_3__T_827_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_6_3__T_315_data; // @[loaf.scala 147:67]
  wire [4:0] AE_6_3__T_315_addr; // @[loaf.scala 147:67]
  wire  AE_6_3__T_315_mask; // @[loaf.scala 147:67]
  wire  AE_6_3__T_315_en; // @[loaf.scala 147:67]
  reg [31:0] AE_6_4 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_52;
  wire [31:0] AE_6_4__T_915_data; // @[loaf.scala 147:67]
  wire [4:0] AE_6_4__T_915_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_6_4__T_321_data; // @[loaf.scala 147:67]
  wire [4:0] AE_6_4__T_321_addr; // @[loaf.scala 147:67]
  wire  AE_6_4__T_321_mask; // @[loaf.scala 147:67]
  wire  AE_6_4__T_321_en; // @[loaf.scala 147:67]
  reg [31:0] AE_6_5 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_53;
  wire [31:0] AE_6_5__T_1003_data; // @[loaf.scala 147:67]
  wire [4:0] AE_6_5__T_1003_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_6_5__T_327_data; // @[loaf.scala 147:67]
  wire [4:0] AE_6_5__T_327_addr; // @[loaf.scala 147:67]
  wire  AE_6_5__T_327_mask; // @[loaf.scala 147:67]
  wire  AE_6_5__T_327_en; // @[loaf.scala 147:67]
  reg [31:0] AE_6_6 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_54;
  wire [31:0] AE_6_6__T_1091_data; // @[loaf.scala 147:67]
  wire [4:0] AE_6_6__T_1091_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_6_6__T_333_data; // @[loaf.scala 147:67]
  wire [4:0] AE_6_6__T_333_addr; // @[loaf.scala 147:67]
  wire  AE_6_6__T_333_mask; // @[loaf.scala 147:67]
  wire  AE_6_6__T_333_en; // @[loaf.scala 147:67]
  reg [31:0] AE_6_7 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_55;
  wire [31:0] AE_6_7__T_1179_data; // @[loaf.scala 147:67]
  wire [4:0] AE_6_7__T_1179_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_6_7__T_339_data; // @[loaf.scala 147:67]
  wire [4:0] AE_6_7__T_339_addr; // @[loaf.scala 147:67]
  wire  AE_6_7__T_339_mask; // @[loaf.scala 147:67]
  wire  AE_6_7__T_339_en; // @[loaf.scala 147:67]
  reg [31:0] AE_7_0 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_56;
  wire [31:0] AE_7_0__T_574_data; // @[loaf.scala 147:67]
  wire [4:0] AE_7_0__T_574_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_7_0__T_345_data; // @[loaf.scala 147:67]
  wire [4:0] AE_7_0__T_345_addr; // @[loaf.scala 147:67]
  wire  AE_7_0__T_345_mask; // @[loaf.scala 147:67]
  wire  AE_7_0__T_345_en; // @[loaf.scala 147:67]
  reg [31:0] AE_7_1 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_57;
  wire [31:0] AE_7_1__T_662_data; // @[loaf.scala 147:67]
  wire [4:0] AE_7_1__T_662_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_7_1__T_351_data; // @[loaf.scala 147:67]
  wire [4:0] AE_7_1__T_351_addr; // @[loaf.scala 147:67]
  wire  AE_7_1__T_351_mask; // @[loaf.scala 147:67]
  wire  AE_7_1__T_351_en; // @[loaf.scala 147:67]
  reg [31:0] AE_7_2 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_58;
  wire [31:0] AE_7_2__T_750_data; // @[loaf.scala 147:67]
  wire [4:0] AE_7_2__T_750_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_7_2__T_357_data; // @[loaf.scala 147:67]
  wire [4:0] AE_7_2__T_357_addr; // @[loaf.scala 147:67]
  wire  AE_7_2__T_357_mask; // @[loaf.scala 147:67]
  wire  AE_7_2__T_357_en; // @[loaf.scala 147:67]
  reg [31:0] AE_7_3 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_59;
  wire [31:0] AE_7_3__T_838_data; // @[loaf.scala 147:67]
  wire [4:0] AE_7_3__T_838_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_7_3__T_363_data; // @[loaf.scala 147:67]
  wire [4:0] AE_7_3__T_363_addr; // @[loaf.scala 147:67]
  wire  AE_7_3__T_363_mask; // @[loaf.scala 147:67]
  wire  AE_7_3__T_363_en; // @[loaf.scala 147:67]
  reg [31:0] AE_7_4 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_60;
  wire [31:0] AE_7_4__T_926_data; // @[loaf.scala 147:67]
  wire [4:0] AE_7_4__T_926_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_7_4__T_369_data; // @[loaf.scala 147:67]
  wire [4:0] AE_7_4__T_369_addr; // @[loaf.scala 147:67]
  wire  AE_7_4__T_369_mask; // @[loaf.scala 147:67]
  wire  AE_7_4__T_369_en; // @[loaf.scala 147:67]
  reg [31:0] AE_7_5 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_61;
  wire [31:0] AE_7_5__T_1014_data; // @[loaf.scala 147:67]
  wire [4:0] AE_7_5__T_1014_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_7_5__T_375_data; // @[loaf.scala 147:67]
  wire [4:0] AE_7_5__T_375_addr; // @[loaf.scala 147:67]
  wire  AE_7_5__T_375_mask; // @[loaf.scala 147:67]
  wire  AE_7_5__T_375_en; // @[loaf.scala 147:67]
  reg [31:0] AE_7_6 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_62;
  wire [31:0] AE_7_6__T_1102_data; // @[loaf.scala 147:67]
  wire [4:0] AE_7_6__T_1102_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_7_6__T_381_data; // @[loaf.scala 147:67]
  wire [4:0] AE_7_6__T_381_addr; // @[loaf.scala 147:67]
  wire  AE_7_6__T_381_mask; // @[loaf.scala 147:67]
  wire  AE_7_6__T_381_en; // @[loaf.scala 147:67]
  reg [31:0] AE_7_7 [0:31]; // @[loaf.scala 147:67]
  reg [31:0] _RAND_63;
  wire [31:0] AE_7_7__T_1190_data; // @[loaf.scala 147:67]
  wire [4:0] AE_7_7__T_1190_addr; // @[loaf.scala 147:67]
  wire [31:0] AE_7_7__T_387_data; // @[loaf.scala 147:67]
  wire [4:0] AE_7_7__T_387_addr; // @[loaf.scala 147:67]
  wire  AE_7_7__T_387_mask; // @[loaf.scala 147:67]
  wire  AE_7_7__T_387_en; // @[loaf.scala 147:67]
  reg [8:0] islice; // @[loaf.scala 108:23]
  reg [31:0] _RAND_64;
  reg  done; // @[loaf.scala 109:21]
  reg [31:0] _RAND_65;
  reg  phase; // @[loaf.scala 111:22]
  reg [31:0] _RAND_66;
  reg [15:0] offCLs_0_0; // @[loaf.scala 113:19]
  reg [31:0] _RAND_67;
  reg [15:0] offCLs_0_1; // @[loaf.scala 113:19]
  reg [31:0] _RAND_68;
  reg [15:0] offCLs_0_2; // @[loaf.scala 113:19]
  reg [31:0] _RAND_69;
  reg [15:0] offCLs_0_3; // @[loaf.scala 113:19]
  reg [31:0] _RAND_70;
  reg [15:0] offCLs_0_4; // @[loaf.scala 113:19]
  reg [31:0] _RAND_71;
  reg [15:0] offCLs_0_5; // @[loaf.scala 113:19]
  reg [31:0] _RAND_72;
  reg [15:0] offCLs_0_6; // @[loaf.scala 113:19]
  reg [31:0] _RAND_73;
  reg [15:0] offCLs_0_7; // @[loaf.scala 113:19]
  reg [31:0] _RAND_74;
  reg [15:0] offCLs_1_0; // @[loaf.scala 113:19]
  reg [31:0] _RAND_75;
  reg [15:0] offCLs_1_1; // @[loaf.scala 113:19]
  reg [31:0] _RAND_76;
  reg [15:0] offCLs_1_2; // @[loaf.scala 113:19]
  reg [31:0] _RAND_77;
  reg [15:0] offCLs_1_3; // @[loaf.scala 113:19]
  reg [31:0] _RAND_78;
  reg [15:0] offCLs_1_4; // @[loaf.scala 113:19]
  reg [31:0] _RAND_79;
  reg [15:0] offCLs_1_5; // @[loaf.scala 113:19]
  reg [31:0] _RAND_80;
  reg [15:0] offCLs_1_6; // @[loaf.scala 113:19]
  reg [31:0] _RAND_81;
  reg [15:0] offCLs_1_7; // @[loaf.scala 113:19]
  reg [31:0] _RAND_82;
  reg [15:0] offCLs_2_0; // @[loaf.scala 113:19]
  reg [31:0] _RAND_83;
  reg [15:0] offCLs_2_1; // @[loaf.scala 113:19]
  reg [31:0] _RAND_84;
  reg [15:0] offCLs_2_2; // @[loaf.scala 113:19]
  reg [31:0] _RAND_85;
  reg [15:0] offCLs_2_3; // @[loaf.scala 113:19]
  reg [31:0] _RAND_86;
  reg [15:0] offCLs_2_4; // @[loaf.scala 113:19]
  reg [31:0] _RAND_87;
  reg [15:0] offCLs_2_5; // @[loaf.scala 113:19]
  reg [31:0] _RAND_88;
  reg [15:0] offCLs_2_6; // @[loaf.scala 113:19]
  reg [31:0] _RAND_89;
  reg [15:0] offCLs_2_7; // @[loaf.scala 113:19]
  reg [31:0] _RAND_90;
  reg [15:0] offCLs_3_0; // @[loaf.scala 113:19]
  reg [31:0] _RAND_91;
  reg [15:0] offCLs_3_1; // @[loaf.scala 113:19]
  reg [31:0] _RAND_92;
  reg [15:0] offCLs_3_2; // @[loaf.scala 113:19]
  reg [31:0] _RAND_93;
  reg [15:0] offCLs_3_3; // @[loaf.scala 113:19]
  reg [31:0] _RAND_94;
  reg [15:0] offCLs_3_4; // @[loaf.scala 113:19]
  reg [31:0] _RAND_95;
  reg [15:0] offCLs_3_5; // @[loaf.scala 113:19]
  reg [31:0] _RAND_96;
  reg [15:0] offCLs_3_6; // @[loaf.scala 113:19]
  reg [31:0] _RAND_97;
  reg [15:0] offCLs_3_7; // @[loaf.scala 113:19]
  reg [31:0] _RAND_98;
  reg [15:0] o1_0; // @[loaf.scala 115:15]
  reg [31:0] _RAND_99;
  reg [15:0] o1_1; // @[loaf.scala 115:15]
  reg [31:0] _RAND_100;
  reg [15:0] o1_2; // @[loaf.scala 115:15]
  reg [31:0] _RAND_101;
  reg [15:0] o1_3; // @[loaf.scala 115:15]
  reg [31:0] _RAND_102;
  reg [15:0] o1_4; // @[loaf.scala 115:15]
  reg [31:0] _RAND_103;
  reg [15:0] o1_5; // @[loaf.scala 115:15]
  reg [31:0] _RAND_104;
  reg [15:0] o1_6; // @[loaf.scala 115:15]
  reg [31:0] _RAND_105;
  reg [15:0] o1_7; // @[loaf.scala 115:15]
  reg [31:0] _RAND_106;
  reg [15:0] o2_0; // @[loaf.scala 116:15]
  reg [31:0] _RAND_107;
  reg [15:0] o2_1; // @[loaf.scala 116:15]
  reg [31:0] _RAND_108;
  reg [15:0] o2_2; // @[loaf.scala 116:15]
  reg [31:0] _RAND_109;
  reg [15:0] o2_3; // @[loaf.scala 116:15]
  reg [31:0] _RAND_110;
  reg [15:0] o2_4; // @[loaf.scala 116:15]
  reg [31:0] _RAND_111;
  reg [15:0] o2_5; // @[loaf.scala 116:15]
  reg [31:0] _RAND_112;
  reg [15:0] o2_6; // @[loaf.scala 116:15]
  reg [31:0] _RAND_113;
  reg [15:0] o2_7; // @[loaf.scala 116:15]
  reg [31:0] _RAND_114;
  reg [15:0] mx2_0_0; // @[loaf.scala 117:68]
  reg [31:0] _RAND_115;
  reg [15:0] mx2_0_1; // @[loaf.scala 117:68]
  reg [31:0] _RAND_116;
  reg [15:0] mx2_0_2; // @[loaf.scala 117:68]
  reg [31:0] _RAND_117;
  reg [15:0] mx2_0_3; // @[loaf.scala 117:68]
  reg [31:0] _RAND_118;
  reg [15:0] mx2_0_4; // @[loaf.scala 117:68]
  reg [31:0] _RAND_119;
  reg [15:0] mx2_0_5; // @[loaf.scala 117:68]
  reg [31:0] _RAND_120;
  reg [15:0] mx2_0_6; // @[loaf.scala 117:68]
  reg [31:0] _RAND_121;
  reg [15:0] mx2_0_7; // @[loaf.scala 117:68]
  reg [31:0] _RAND_122;
  reg [15:0] mx2_1_0; // @[loaf.scala 117:68]
  reg [31:0] _RAND_123;
  reg [15:0] mx2_1_1; // @[loaf.scala 117:68]
  reg [31:0] _RAND_124;
  reg [15:0] mx2_1_2; // @[loaf.scala 117:68]
  reg [31:0] _RAND_125;
  reg [15:0] mx2_1_3; // @[loaf.scala 117:68]
  reg [31:0] _RAND_126;
  reg [15:0] mx2_1_4; // @[loaf.scala 117:68]
  reg [31:0] _RAND_127;
  reg [15:0] mx2_1_5; // @[loaf.scala 117:68]
  reg [31:0] _RAND_128;
  reg [15:0] mx2_1_6; // @[loaf.scala 117:68]
  reg [31:0] _RAND_129;
  reg [15:0] mx2_1_7; // @[loaf.scala 117:68]
  reg [31:0] _RAND_130;
  reg [15:0] mx2_2_0; // @[loaf.scala 117:68]
  reg [31:0] _RAND_131;
  reg [15:0] mx2_2_1; // @[loaf.scala 117:68]
  reg [31:0] _RAND_132;
  reg [15:0] mx2_2_2; // @[loaf.scala 117:68]
  reg [31:0] _RAND_133;
  reg [15:0] mx2_2_3; // @[loaf.scala 117:68]
  reg [31:0] _RAND_134;
  reg [15:0] mx2_2_4; // @[loaf.scala 117:68]
  reg [31:0] _RAND_135;
  reg [15:0] mx2_2_5; // @[loaf.scala 117:68]
  reg [31:0] _RAND_136;
  reg [15:0] mx2_2_6; // @[loaf.scala 117:68]
  reg [31:0] _RAND_137;
  reg [15:0] mx2_2_7; // @[loaf.scala 117:68]
  reg [31:0] _RAND_138;
  reg [15:0] mx2_3_0; // @[loaf.scala 117:68]
  reg [31:0] _RAND_139;
  reg [15:0] mx2_3_1; // @[loaf.scala 117:68]
  reg [31:0] _RAND_140;
  reg [15:0] mx2_3_2; // @[loaf.scala 117:68]
  reg [31:0] _RAND_141;
  reg [15:0] mx2_3_3; // @[loaf.scala 117:68]
  reg [31:0] _RAND_142;
  reg [15:0] mx2_3_4; // @[loaf.scala 117:68]
  reg [31:0] _RAND_143;
  reg [15:0] mx2_3_5; // @[loaf.scala 117:68]
  reg [31:0] _RAND_144;
  reg [15:0] mx2_3_6; // @[loaf.scala 117:68]
  reg [31:0] _RAND_145;
  reg [15:0] mx2_3_7; // @[loaf.scala 117:68]
  reg [31:0] _RAND_146;
  reg [15:0] mx2_4_0; // @[loaf.scala 117:68]
  reg [31:0] _RAND_147;
  reg [15:0] mx2_4_1; // @[loaf.scala 117:68]
  reg [31:0] _RAND_148;
  reg [15:0] mx2_4_2; // @[loaf.scala 117:68]
  reg [31:0] _RAND_149;
  reg [15:0] mx2_4_3; // @[loaf.scala 117:68]
  reg [31:0] _RAND_150;
  reg [15:0] mx2_4_4; // @[loaf.scala 117:68]
  reg [31:0] _RAND_151;
  reg [15:0] mx2_4_5; // @[loaf.scala 117:68]
  reg [31:0] _RAND_152;
  reg [15:0] mx2_4_6; // @[loaf.scala 117:68]
  reg [31:0] _RAND_153;
  reg [15:0] mx2_4_7; // @[loaf.scala 117:68]
  reg [31:0] _RAND_154;
  reg [15:0] mx2_5_0; // @[loaf.scala 117:68]
  reg [31:0] _RAND_155;
  reg [15:0] mx2_5_1; // @[loaf.scala 117:68]
  reg [31:0] _RAND_156;
  reg [15:0] mx2_5_2; // @[loaf.scala 117:68]
  reg [31:0] _RAND_157;
  reg [15:0] mx2_5_3; // @[loaf.scala 117:68]
  reg [31:0] _RAND_158;
  reg [15:0] mx2_5_4; // @[loaf.scala 117:68]
  reg [31:0] _RAND_159;
  reg [15:0] mx2_5_5; // @[loaf.scala 117:68]
  reg [31:0] _RAND_160;
  reg [15:0] mx2_5_6; // @[loaf.scala 117:68]
  reg [31:0] _RAND_161;
  reg [15:0] mx2_5_7; // @[loaf.scala 117:68]
  reg [31:0] _RAND_162;
  reg [15:0] mx2_6_0; // @[loaf.scala 117:68]
  reg [31:0] _RAND_163;
  reg [15:0] mx2_6_1; // @[loaf.scala 117:68]
  reg [31:0] _RAND_164;
  reg [15:0] mx2_6_2; // @[loaf.scala 117:68]
  reg [31:0] _RAND_165;
  reg [15:0] mx2_6_3; // @[loaf.scala 117:68]
  reg [31:0] _RAND_166;
  reg [15:0] mx2_6_4; // @[loaf.scala 117:68]
  reg [31:0] _RAND_167;
  reg [15:0] mx2_6_5; // @[loaf.scala 117:68]
  reg [31:0] _RAND_168;
  reg [15:0] mx2_6_6; // @[loaf.scala 117:68]
  reg [31:0] _RAND_169;
  reg [15:0] mx2_6_7; // @[loaf.scala 117:68]
  reg [31:0] _RAND_170;
  reg [15:0] mx2_7_0; // @[loaf.scala 117:68]
  reg [31:0] _RAND_171;
  reg [15:0] mx2_7_1; // @[loaf.scala 117:68]
  reg [31:0] _RAND_172;
  reg [15:0] mx2_7_2; // @[loaf.scala 117:68]
  reg [31:0] _RAND_173;
  reg [15:0] mx2_7_3; // @[loaf.scala 117:68]
  reg [31:0] _RAND_174;
  reg [15:0] mx2_7_4; // @[loaf.scala 117:68]
  reg [31:0] _RAND_175;
  reg [15:0] mx2_7_5; // @[loaf.scala 117:68]
  reg [31:0] _RAND_176;
  reg [15:0] mx2_7_6; // @[loaf.scala 117:68]
  reg [31:0] _RAND_177;
  reg [15:0] mx2_7_7; // @[loaf.scala 117:68]
  reg [31:0] _RAND_178;
  reg [15:0] ab2_0_0; // @[loaf.scala 118:68]
  reg [31:0] _RAND_179;
  reg [15:0] ab2_0_1; // @[loaf.scala 118:68]
  reg [31:0] _RAND_180;
  reg [15:0] ab2_0_2; // @[loaf.scala 118:68]
  reg [31:0] _RAND_181;
  reg [15:0] ab2_0_3; // @[loaf.scala 118:68]
  reg [31:0] _RAND_182;
  reg [15:0] ab2_0_4; // @[loaf.scala 118:68]
  reg [31:0] _RAND_183;
  reg [15:0] ab2_0_5; // @[loaf.scala 118:68]
  reg [31:0] _RAND_184;
  reg [15:0] ab2_0_6; // @[loaf.scala 118:68]
  reg [31:0] _RAND_185;
  reg [15:0] ab2_0_7; // @[loaf.scala 118:68]
  reg [31:0] _RAND_186;
  reg [15:0] ab2_1_0; // @[loaf.scala 118:68]
  reg [31:0] _RAND_187;
  reg [15:0] ab2_1_1; // @[loaf.scala 118:68]
  reg [31:0] _RAND_188;
  reg [15:0] ab2_1_2; // @[loaf.scala 118:68]
  reg [31:0] _RAND_189;
  reg [15:0] ab2_1_3; // @[loaf.scala 118:68]
  reg [31:0] _RAND_190;
  reg [15:0] ab2_1_4; // @[loaf.scala 118:68]
  reg [31:0] _RAND_191;
  reg [15:0] ab2_1_5; // @[loaf.scala 118:68]
  reg [31:0] _RAND_192;
  reg [15:0] ab2_1_6; // @[loaf.scala 118:68]
  reg [31:0] _RAND_193;
  reg [15:0] ab2_1_7; // @[loaf.scala 118:68]
  reg [31:0] _RAND_194;
  reg [15:0] ab2_2_0; // @[loaf.scala 118:68]
  reg [31:0] _RAND_195;
  reg [15:0] ab2_2_1; // @[loaf.scala 118:68]
  reg [31:0] _RAND_196;
  reg [15:0] ab2_2_2; // @[loaf.scala 118:68]
  reg [31:0] _RAND_197;
  reg [15:0] ab2_2_3; // @[loaf.scala 118:68]
  reg [31:0] _RAND_198;
  reg [15:0] ab2_2_4; // @[loaf.scala 118:68]
  reg [31:0] _RAND_199;
  reg [15:0] ab2_2_5; // @[loaf.scala 118:68]
  reg [31:0] _RAND_200;
  reg [15:0] ab2_2_6; // @[loaf.scala 118:68]
  reg [31:0] _RAND_201;
  reg [15:0] ab2_2_7; // @[loaf.scala 118:68]
  reg [31:0] _RAND_202;
  reg [15:0] ab2_3_0; // @[loaf.scala 118:68]
  reg [31:0] _RAND_203;
  reg [15:0] ab2_3_1; // @[loaf.scala 118:68]
  reg [31:0] _RAND_204;
  reg [15:0] ab2_3_2; // @[loaf.scala 118:68]
  reg [31:0] _RAND_205;
  reg [15:0] ab2_3_3; // @[loaf.scala 118:68]
  reg [31:0] _RAND_206;
  reg [15:0] ab2_3_4; // @[loaf.scala 118:68]
  reg [31:0] _RAND_207;
  reg [15:0] ab2_3_5; // @[loaf.scala 118:68]
  reg [31:0] _RAND_208;
  reg [15:0] ab2_3_6; // @[loaf.scala 118:68]
  reg [31:0] _RAND_209;
  reg [15:0] ab2_3_7; // @[loaf.scala 118:68]
  reg [31:0] _RAND_210;
  reg [15:0] ab2_4_0; // @[loaf.scala 118:68]
  reg [31:0] _RAND_211;
  reg [15:0] ab2_4_1; // @[loaf.scala 118:68]
  reg [31:0] _RAND_212;
  reg [15:0] ab2_4_2; // @[loaf.scala 118:68]
  reg [31:0] _RAND_213;
  reg [15:0] ab2_4_3; // @[loaf.scala 118:68]
  reg [31:0] _RAND_214;
  reg [15:0] ab2_4_4; // @[loaf.scala 118:68]
  reg [31:0] _RAND_215;
  reg [15:0] ab2_4_5; // @[loaf.scala 118:68]
  reg [31:0] _RAND_216;
  reg [15:0] ab2_4_6; // @[loaf.scala 118:68]
  reg [31:0] _RAND_217;
  reg [15:0] ab2_4_7; // @[loaf.scala 118:68]
  reg [31:0] _RAND_218;
  reg [15:0] ab2_5_0; // @[loaf.scala 118:68]
  reg [31:0] _RAND_219;
  reg [15:0] ab2_5_1; // @[loaf.scala 118:68]
  reg [31:0] _RAND_220;
  reg [15:0] ab2_5_2; // @[loaf.scala 118:68]
  reg [31:0] _RAND_221;
  reg [15:0] ab2_5_3; // @[loaf.scala 118:68]
  reg [31:0] _RAND_222;
  reg [15:0] ab2_5_4; // @[loaf.scala 118:68]
  reg [31:0] _RAND_223;
  reg [15:0] ab2_5_5; // @[loaf.scala 118:68]
  reg [31:0] _RAND_224;
  reg [15:0] ab2_5_6; // @[loaf.scala 118:68]
  reg [31:0] _RAND_225;
  reg [15:0] ab2_5_7; // @[loaf.scala 118:68]
  reg [31:0] _RAND_226;
  reg [15:0] ab2_6_0; // @[loaf.scala 118:68]
  reg [31:0] _RAND_227;
  reg [15:0] ab2_6_1; // @[loaf.scala 118:68]
  reg [31:0] _RAND_228;
  reg [15:0] ab2_6_2; // @[loaf.scala 118:68]
  reg [31:0] _RAND_229;
  reg [15:0] ab2_6_3; // @[loaf.scala 118:68]
  reg [31:0] _RAND_230;
  reg [15:0] ab2_6_4; // @[loaf.scala 118:68]
  reg [31:0] _RAND_231;
  reg [15:0] ab2_6_5; // @[loaf.scala 118:68]
  reg [31:0] _RAND_232;
  reg [15:0] ab2_6_6; // @[loaf.scala 118:68]
  reg [31:0] _RAND_233;
  reg [15:0] ab2_6_7; // @[loaf.scala 118:68]
  reg [31:0] _RAND_234;
  reg [15:0] ab2_7_0; // @[loaf.scala 118:68]
  reg [31:0] _RAND_235;
  reg [15:0] ab2_7_1; // @[loaf.scala 118:68]
  reg [31:0] _RAND_236;
  reg [15:0] ab2_7_2; // @[loaf.scala 118:68]
  reg [31:0] _RAND_237;
  reg [15:0] ab2_7_3; // @[loaf.scala 118:68]
  reg [31:0] _RAND_238;
  reg [15:0] ab2_7_4; // @[loaf.scala 118:68]
  reg [31:0] _RAND_239;
  reg [15:0] ab2_7_5; // @[loaf.scala 118:68]
  reg [31:0] _RAND_240;
  reg [15:0] ab2_7_6; // @[loaf.scala 118:68]
  reg [31:0] _RAND_241;
  reg [15:0] ab2_7_7; // @[loaf.scala 118:68]
  reg [31:0] _RAND_242;
  reg [15:0] tm8_0_0; // @[loaf.scala 122:82]
  reg [31:0] _RAND_243;
  reg [15:0] tm8_0_1; // @[loaf.scala 122:82]
  reg [31:0] _RAND_244;
  reg [15:0] tm8_0_2; // @[loaf.scala 122:82]
  reg [31:0] _RAND_245;
  reg [15:0] tm8_0_3; // @[loaf.scala 122:82]
  reg [31:0] _RAND_246;
  reg [15:0] tm8_0_4; // @[loaf.scala 122:82]
  reg [31:0] _RAND_247;
  reg [15:0] tm8_0_5; // @[loaf.scala 122:82]
  reg [31:0] _RAND_248;
  reg [15:0] tm8_0_6; // @[loaf.scala 122:82]
  reg [31:0] _RAND_249;
  reg [15:0] tm8_0_7; // @[loaf.scala 122:82]
  reg [31:0] _RAND_250;
  reg [15:0] tm8_1_0; // @[loaf.scala 122:82]
  reg [31:0] _RAND_251;
  reg [15:0] tm8_1_1; // @[loaf.scala 122:82]
  reg [31:0] _RAND_252;
  reg [15:0] tm8_1_2; // @[loaf.scala 122:82]
  reg [31:0] _RAND_253;
  reg [15:0] tm8_1_3; // @[loaf.scala 122:82]
  reg [31:0] _RAND_254;
  reg [15:0] tm8_1_4; // @[loaf.scala 122:82]
  reg [31:0] _RAND_255;
  reg [15:0] tm8_1_5; // @[loaf.scala 122:82]
  reg [31:0] _RAND_256;
  reg [15:0] tm8_1_6; // @[loaf.scala 122:82]
  reg [31:0] _RAND_257;
  reg [15:0] tm8_1_7; // @[loaf.scala 122:82]
  reg [31:0] _RAND_258;
  reg [15:0] tm8_2_0; // @[loaf.scala 122:82]
  reg [31:0] _RAND_259;
  reg [15:0] tm8_2_1; // @[loaf.scala 122:82]
  reg [31:0] _RAND_260;
  reg [15:0] tm8_2_2; // @[loaf.scala 122:82]
  reg [31:0] _RAND_261;
  reg [15:0] tm8_2_3; // @[loaf.scala 122:82]
  reg [31:0] _RAND_262;
  reg [15:0] tm8_2_4; // @[loaf.scala 122:82]
  reg [31:0] _RAND_263;
  reg [15:0] tm8_2_5; // @[loaf.scala 122:82]
  reg [31:0] _RAND_264;
  reg [15:0] tm8_2_6; // @[loaf.scala 122:82]
  reg [31:0] _RAND_265;
  reg [15:0] tm8_2_7; // @[loaf.scala 122:82]
  reg [31:0] _RAND_266;
  reg [15:0] tm8_3_0; // @[loaf.scala 122:82]
  reg [31:0] _RAND_267;
  reg [15:0] tm8_3_1; // @[loaf.scala 122:82]
  reg [31:0] _RAND_268;
  reg [15:0] tm8_3_2; // @[loaf.scala 122:82]
  reg [31:0] _RAND_269;
  reg [15:0] tm8_3_3; // @[loaf.scala 122:82]
  reg [31:0] _RAND_270;
  reg [15:0] tm8_3_4; // @[loaf.scala 122:82]
  reg [31:0] _RAND_271;
  reg [15:0] tm8_3_5; // @[loaf.scala 122:82]
  reg [31:0] _RAND_272;
  reg [15:0] tm8_3_6; // @[loaf.scala 122:82]
  reg [31:0] _RAND_273;
  reg [15:0] tm8_3_7; // @[loaf.scala 122:82]
  reg [31:0] _RAND_274;
  reg [15:0] tm9_0_0; // @[loaf.scala 123:82]
  reg [31:0] _RAND_275;
  reg [15:0] tm9_0_1; // @[loaf.scala 123:82]
  reg [31:0] _RAND_276;
  reg [15:0] tm9_0_2; // @[loaf.scala 123:82]
  reg [31:0] _RAND_277;
  reg [15:0] tm9_0_3; // @[loaf.scala 123:82]
  reg [31:0] _RAND_278;
  reg [15:0] tm9_0_4; // @[loaf.scala 123:82]
  reg [31:0] _RAND_279;
  reg [15:0] tm9_0_5; // @[loaf.scala 123:82]
  reg [31:0] _RAND_280;
  reg [15:0] tm9_0_6; // @[loaf.scala 123:82]
  reg [31:0] _RAND_281;
  reg [15:0] tm9_0_7; // @[loaf.scala 123:82]
  reg [31:0] _RAND_282;
  reg [15:0] tm9_1_0; // @[loaf.scala 123:82]
  reg [31:0] _RAND_283;
  reg [15:0] tm9_1_1; // @[loaf.scala 123:82]
  reg [31:0] _RAND_284;
  reg [15:0] tm9_1_2; // @[loaf.scala 123:82]
  reg [31:0] _RAND_285;
  reg [15:0] tm9_1_3; // @[loaf.scala 123:82]
  reg [31:0] _RAND_286;
  reg [15:0] tm9_1_4; // @[loaf.scala 123:82]
  reg [31:0] _RAND_287;
  reg [15:0] tm9_1_5; // @[loaf.scala 123:82]
  reg [31:0] _RAND_288;
  reg [15:0] tm9_1_6; // @[loaf.scala 123:82]
  reg [31:0] _RAND_289;
  reg [15:0] tm9_1_7; // @[loaf.scala 123:82]
  reg [31:0] _RAND_290;
  reg [15:0] tma_0_0; // @[loaf.scala 124:82]
  reg [31:0] _RAND_291;
  reg [15:0] tma_0_1; // @[loaf.scala 124:82]
  reg [31:0] _RAND_292;
  reg [15:0] tma_0_2; // @[loaf.scala 124:82]
  reg [31:0] _RAND_293;
  reg [15:0] tma_0_3; // @[loaf.scala 124:82]
  reg [31:0] _RAND_294;
  reg [15:0] tma_0_4; // @[loaf.scala 124:82]
  reg [31:0] _RAND_295;
  reg [15:0] tma_0_5; // @[loaf.scala 124:82]
  reg [31:0] _RAND_296;
  reg [15:0] tma_0_6; // @[loaf.scala 124:82]
  reg [31:0] _RAND_297;
  reg [15:0] tma_0_7; // @[loaf.scala 124:82]
  reg [31:0] _RAND_298;
  reg [15:0] tmb_0_0; // @[loaf.scala 125:82]
  reg [31:0] _RAND_299;
  reg [15:0] tmb_0_1; // @[loaf.scala 125:82]
  reg [31:0] _RAND_300;
  reg [15:0] tmb_0_2; // @[loaf.scala 125:82]
  reg [31:0] _RAND_301;
  reg [15:0] tmb_0_3; // @[loaf.scala 125:82]
  reg [31:0] _RAND_302;
  reg [15:0] tmb_0_4; // @[loaf.scala 125:82]
  reg [31:0] _RAND_303;
  reg [15:0] tmb_0_5; // @[loaf.scala 125:82]
  reg [31:0] _RAND_304;
  reg [15:0] tmb_0_6; // @[loaf.scala 125:82]
  reg [31:0] _RAND_305;
  reg [15:0] tmb_0_7; // @[loaf.scala 125:82]
  reg [31:0] _RAND_306;
  reg [15:0] tmc_0_0; // @[loaf.scala 126:82]
  reg [31:0] _RAND_307;
  reg [15:0] tmc_0_1; // @[loaf.scala 126:82]
  reg [31:0] _RAND_308;
  reg [15:0] tmc_0_2; // @[loaf.scala 126:82]
  reg [31:0] _RAND_309;
  reg [15:0] tmc_0_3; // @[loaf.scala 126:82]
  reg [31:0] _RAND_310;
  reg [15:0] tmc_0_4; // @[loaf.scala 126:82]
  reg [31:0] _RAND_311;
  reg [15:0] tmc_0_5; // @[loaf.scala 126:82]
  reg [31:0] _RAND_312;
  reg [15:0] tmc_0_6; // @[loaf.scala 126:82]
  reg [31:0] _RAND_313;
  reg [15:0] tmc_0_7; // @[loaf.scala 126:82]
  reg [31:0] _RAND_314;
  reg [15:0] best_0; // @[loaf.scala 128:17]
  reg [31:0] _RAND_315;
  reg [15:0] best_1; // @[loaf.scala 128:17]
  reg [31:0] _RAND_316;
  reg [15:0] best_2; // @[loaf.scala 128:17]
  reg [31:0] _RAND_317;
  reg [15:0] best_3; // @[loaf.scala 128:17]
  reg [31:0] _RAND_318;
  reg [15:0] best_4; // @[loaf.scala 128:17]
  reg [31:0] _RAND_319;
  reg [15:0] best_5; // @[loaf.scala 128:17]
  reg [31:0] _RAND_320;
  reg [15:0] best_6; // @[loaf.scala 128:17]
  reg [31:0] _RAND_321;
  reg [15:0] best_7; // @[loaf.scala 128:17]
  reg [31:0] _RAND_322;
  reg [15:0] bestBufe_0; // @[loaf.scala 129:21]
  reg [31:0] _RAND_323;
  reg [15:0] bestBufe_1; // @[loaf.scala 129:21]
  reg [31:0] _RAND_324;
  reg [15:0] bestBufe_2; // @[loaf.scala 129:21]
  reg [31:0] _RAND_325;
  reg [15:0] bestBufe_3; // @[loaf.scala 129:21]
  reg [31:0] _RAND_326;
  reg [15:0] bestBufe_4; // @[loaf.scala 129:21]
  reg [31:0] _RAND_327;
  reg [15:0] bestBufe_5; // @[loaf.scala 129:21]
  reg [31:0] _RAND_328;
  reg [15:0] bestBufe_6; // @[loaf.scala 129:21]
  reg [31:0] _RAND_329;
  reg [15:0] bestBufe_7; // @[loaf.scala 129:21]
  reg [31:0] _RAND_330;
  reg [1:0] r; // @[loaf.scala 131:18]
  reg [31:0] _RAND_331;
  reg [1:0] c; // @[loaf.scala 132:18]
  reg [31:0] _RAND_332;
  reg [15:0] BFbuf_e; // @[loaf.scala 134:18]
  reg [31:0] _RAND_333;
  reg [15:0] BFbuf_a; // @[loaf.scala 134:18]
  reg [31:0] _RAND_334;
  reg [4:0] load_i; // @[loaf.scala 136:23]
  reg [31:0] _RAND_335;
  reg [4:0] load_j; // @[loaf.scala 137:23]
  reg [31:0] _RAND_336;
  reg  doneLoading; // @[loaf.scala 138:28]
  reg [31:0] _RAND_337;
  reg  lastLoad; // @[loaf.scala 139:25]
  reg [31:0] _RAND_338;
  reg [2:0] prev_lo_i; // @[loaf.scala 141:22]
  reg [31:0] _RAND_339;
  reg [2:0] prev_lo_j; // @[loaf.scala 142:22]
  reg [31:0] _RAND_340;
  reg [4:0] prev_idx; // @[loaf.scala 143:22]
  reg [31:0] _RAND_341;
  reg [15:0] slcBuf_e; // @[loaf.scala 144:19]
  reg [31:0] _RAND_342;
  reg [15:0] slcBuf_a; // @[loaf.scala 144:19]
  reg [31:0] _RAND_343;
  reg  slcValid; // @[loaf.scala 145:25]
  reg [31:0] _RAND_344;
  reg [15:0] AEbuf_0_0_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_345;
  reg [15:0] AEbuf_0_0_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_346;
  reg [15:0] AEbuf_0_1_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_347;
  reg [15:0] AEbuf_0_1_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_348;
  reg [15:0] AEbuf_0_2_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_349;
  reg [15:0] AEbuf_0_2_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_350;
  reg [15:0] AEbuf_0_3_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_351;
  reg [15:0] AEbuf_0_3_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_352;
  reg [15:0] AEbuf_0_4_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_353;
  reg [15:0] AEbuf_0_4_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_354;
  reg [15:0] AEbuf_0_5_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_355;
  reg [15:0] AEbuf_0_5_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_356;
  reg [15:0] AEbuf_0_6_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_357;
  reg [15:0] AEbuf_0_6_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_358;
  reg [15:0] AEbuf_0_7_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_359;
  reg [15:0] AEbuf_0_7_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_360;
  reg [15:0] AEbuf_1_0_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_361;
  reg [15:0] AEbuf_1_0_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_362;
  reg [15:0] AEbuf_1_1_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_363;
  reg [15:0] AEbuf_1_1_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_364;
  reg [15:0] AEbuf_1_2_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_365;
  reg [15:0] AEbuf_1_2_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_366;
  reg [15:0] AEbuf_1_3_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_367;
  reg [15:0] AEbuf_1_3_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_368;
  reg [15:0] AEbuf_1_4_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_369;
  reg [15:0] AEbuf_1_4_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_370;
  reg [15:0] AEbuf_1_5_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_371;
  reg [15:0] AEbuf_1_5_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_372;
  reg [15:0] AEbuf_1_6_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_373;
  reg [15:0] AEbuf_1_6_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_374;
  reg [15:0] AEbuf_1_7_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_375;
  reg [15:0] AEbuf_1_7_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_376;
  reg [15:0] AEbuf_2_0_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_377;
  reg [15:0] AEbuf_2_0_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_378;
  reg [15:0] AEbuf_2_1_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_379;
  reg [15:0] AEbuf_2_1_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_380;
  reg [15:0] AEbuf_2_2_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_381;
  reg [15:0] AEbuf_2_2_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_382;
  reg [15:0] AEbuf_2_3_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_383;
  reg [15:0] AEbuf_2_3_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_384;
  reg [15:0] AEbuf_2_4_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_385;
  reg [15:0] AEbuf_2_4_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_386;
  reg [15:0] AEbuf_2_5_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_387;
  reg [15:0] AEbuf_2_5_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_388;
  reg [15:0] AEbuf_2_6_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_389;
  reg [15:0] AEbuf_2_6_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_390;
  reg [15:0] AEbuf_2_7_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_391;
  reg [15:0] AEbuf_2_7_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_392;
  reg [15:0] AEbuf_3_0_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_393;
  reg [15:0] AEbuf_3_0_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_394;
  reg [15:0] AEbuf_3_1_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_395;
  reg [15:0] AEbuf_3_1_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_396;
  reg [15:0] AEbuf_3_2_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_397;
  reg [15:0] AEbuf_3_2_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_398;
  reg [15:0] AEbuf_3_3_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_399;
  reg [15:0] AEbuf_3_3_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_400;
  reg [15:0] AEbuf_3_4_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_401;
  reg [15:0] AEbuf_3_4_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_402;
  reg [15:0] AEbuf_3_5_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_403;
  reg [15:0] AEbuf_3_5_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_404;
  reg [15:0] AEbuf_3_6_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_405;
  reg [15:0] AEbuf_3_6_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_406;
  reg [15:0] AEbuf_3_7_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_407;
  reg [15:0] AEbuf_3_7_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_408;
  reg [15:0] AEbuf_4_0_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_409;
  reg [15:0] AEbuf_4_0_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_410;
  reg [15:0] AEbuf_4_1_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_411;
  reg [15:0] AEbuf_4_1_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_412;
  reg [15:0] AEbuf_4_2_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_413;
  reg [15:0] AEbuf_4_2_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_414;
  reg [15:0] AEbuf_4_3_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_415;
  reg [15:0] AEbuf_4_3_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_416;
  reg [15:0] AEbuf_4_4_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_417;
  reg [15:0] AEbuf_4_4_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_418;
  reg [15:0] AEbuf_4_5_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_419;
  reg [15:0] AEbuf_4_5_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_420;
  reg [15:0] AEbuf_4_6_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_421;
  reg [15:0] AEbuf_4_6_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_422;
  reg [15:0] AEbuf_4_7_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_423;
  reg [15:0] AEbuf_4_7_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_424;
  reg [15:0] AEbuf_5_0_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_425;
  reg [15:0] AEbuf_5_0_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_426;
  reg [15:0] AEbuf_5_1_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_427;
  reg [15:0] AEbuf_5_1_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_428;
  reg [15:0] AEbuf_5_2_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_429;
  reg [15:0] AEbuf_5_2_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_430;
  reg [15:0] AEbuf_5_3_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_431;
  reg [15:0] AEbuf_5_3_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_432;
  reg [15:0] AEbuf_5_4_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_433;
  reg [15:0] AEbuf_5_4_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_434;
  reg [15:0] AEbuf_5_5_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_435;
  reg [15:0] AEbuf_5_5_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_436;
  reg [15:0] AEbuf_5_6_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_437;
  reg [15:0] AEbuf_5_6_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_438;
  reg [15:0] AEbuf_5_7_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_439;
  reg [15:0] AEbuf_5_7_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_440;
  reg [15:0] AEbuf_6_0_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_441;
  reg [15:0] AEbuf_6_0_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_442;
  reg [15:0] AEbuf_6_1_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_443;
  reg [15:0] AEbuf_6_1_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_444;
  reg [15:0] AEbuf_6_2_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_445;
  reg [15:0] AEbuf_6_2_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_446;
  reg [15:0] AEbuf_6_3_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_447;
  reg [15:0] AEbuf_6_3_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_448;
  reg [15:0] AEbuf_6_4_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_449;
  reg [15:0] AEbuf_6_4_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_450;
  reg [15:0] AEbuf_6_5_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_451;
  reg [15:0] AEbuf_6_5_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_452;
  reg [15:0] AEbuf_6_6_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_453;
  reg [15:0] AEbuf_6_6_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_454;
  reg [15:0] AEbuf_6_7_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_455;
  reg [15:0] AEbuf_6_7_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_456;
  reg [15:0] AEbuf_7_0_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_457;
  reg [15:0] AEbuf_7_0_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_458;
  reg [15:0] AEbuf_7_1_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_459;
  reg [15:0] AEbuf_7_1_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_460;
  reg [15:0] AEbuf_7_2_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_461;
  reg [15:0] AEbuf_7_2_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_462;
  reg [15:0] AEbuf_7_3_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_463;
  reg [15:0] AEbuf_7_3_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_464;
  reg [15:0] AEbuf_7_4_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_465;
  reg [15:0] AEbuf_7_4_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_466;
  reg [15:0] AEbuf_7_5_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_467;
  reg [15:0] AEbuf_7_5_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_468;
  reg [15:0] AEbuf_7_6_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_469;
  reg [15:0] AEbuf_7_6_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_470;
  reg [15:0] AEbuf_7_7_e; // @[loaf.scala 148:70]
  reg [31:0] _RAND_471;
  reg [15:0] AEbuf_7_7_a; // @[loaf.scala 148:70]
  reg [31:0] _RAND_472;
  wire  _T_1; // @[loaf.scala 170:22]
  wire  _T_2; // @[loaf.scala 170:19]
  wire  _T_3; // @[loaf.scala 174:27]
  wire  _T_4; // @[loaf.scala 179:24]
  wire  _T_5; // @[loaf.scala 179:45]
  wire  _T_6; // @[loaf.scala 179:38]
  wire  _T_11; // @[loaf.scala 179:45]
  wire  _T_12; // @[loaf.scala 179:38]
  wire  _T_17; // @[loaf.scala 179:45]
  wire  _T_18; // @[loaf.scala 179:38]
  wire  _T_23; // @[loaf.scala 179:45]
  wire  _T_24; // @[loaf.scala 179:38]
  wire  _T_29; // @[loaf.scala 179:45]
  wire  _T_30; // @[loaf.scala 179:38]
  wire  _T_35; // @[loaf.scala 179:45]
  wire  _T_36; // @[loaf.scala 179:38]
  wire  _T_41; // @[loaf.scala 179:45]
  wire  _T_42; // @[loaf.scala 179:38]
  wire  _T_47; // @[loaf.scala 179:45]
  wire  _T_48; // @[loaf.scala 179:38]
  wire  _T_52; // @[loaf.scala 179:24]
  wire  _T_54; // @[loaf.scala 179:38]
  wire  _T_60; // @[loaf.scala 179:38]
  wire  _T_66; // @[loaf.scala 179:38]
  wire  _T_72; // @[loaf.scala 179:38]
  wire  _T_78; // @[loaf.scala 179:38]
  wire  _T_84; // @[loaf.scala 179:38]
  wire  _T_90; // @[loaf.scala 179:38]
  wire  _T_96; // @[loaf.scala 179:38]
  wire  _T_100; // @[loaf.scala 179:24]
  wire  _T_102; // @[loaf.scala 179:38]
  wire  _T_108; // @[loaf.scala 179:38]
  wire  _T_114; // @[loaf.scala 179:38]
  wire  _T_120; // @[loaf.scala 179:38]
  wire  _T_126; // @[loaf.scala 179:38]
  wire  _T_132; // @[loaf.scala 179:38]
  wire  _T_138; // @[loaf.scala 179:38]
  wire  _T_144; // @[loaf.scala 179:38]
  wire  _T_148; // @[loaf.scala 179:24]
  wire  _T_150; // @[loaf.scala 179:38]
  wire  _T_156; // @[loaf.scala 179:38]
  wire  _T_162; // @[loaf.scala 179:38]
  wire  _T_168; // @[loaf.scala 179:38]
  wire  _T_174; // @[loaf.scala 179:38]
  wire  _T_180; // @[loaf.scala 179:38]
  wire  _T_186; // @[loaf.scala 179:38]
  wire  _T_192; // @[loaf.scala 179:38]
  wire  _T_196; // @[loaf.scala 179:24]
  wire  _T_198; // @[loaf.scala 179:38]
  wire  _T_204; // @[loaf.scala 179:38]
  wire  _T_210; // @[loaf.scala 179:38]
  wire  _T_216; // @[loaf.scala 179:38]
  wire  _T_222; // @[loaf.scala 179:38]
  wire  _T_228; // @[loaf.scala 179:38]
  wire  _T_234; // @[loaf.scala 179:38]
  wire  _T_240; // @[loaf.scala 179:38]
  wire  _T_244; // @[loaf.scala 179:24]
  wire  _T_246; // @[loaf.scala 179:38]
  wire  _T_252; // @[loaf.scala 179:38]
  wire  _T_258; // @[loaf.scala 179:38]
  wire  _T_264; // @[loaf.scala 179:38]
  wire  _T_270; // @[loaf.scala 179:38]
  wire  _T_276; // @[loaf.scala 179:38]
  wire  _T_282; // @[loaf.scala 179:38]
  wire  _T_288; // @[loaf.scala 179:38]
  wire  _T_292; // @[loaf.scala 179:24]
  wire  _T_294; // @[loaf.scala 179:38]
  wire  _T_300; // @[loaf.scala 179:38]
  wire  _T_306; // @[loaf.scala 179:38]
  wire  _T_312; // @[loaf.scala 179:38]
  wire  _T_318; // @[loaf.scala 179:38]
  wire  _T_324; // @[loaf.scala 179:38]
  wire  _T_330; // @[loaf.scala 179:38]
  wire  _T_336; // @[loaf.scala 179:38]
  wire  _T_340; // @[loaf.scala 179:24]
  wire  _T_342; // @[loaf.scala 179:38]
  wire  _T_348; // @[loaf.scala 179:38]
  wire  _T_354; // @[loaf.scala 179:38]
  wire  _T_360; // @[loaf.scala 179:38]
  wire  _T_366; // @[loaf.scala 179:38]
  wire  _T_372; // @[loaf.scala 179:38]
  wire  _T_378; // @[loaf.scala 179:38]
  wire  _T_384; // @[loaf.scala 179:38]
  wire  _GEN_322; // @[loaf.scala 176:26]
  wire  _GEN_327; // @[loaf.scala 176:26]
  wire  _GEN_332; // @[loaf.scala 176:26]
  wire  _GEN_337; // @[loaf.scala 176:26]
  wire  _GEN_342; // @[loaf.scala 176:26]
  wire  _GEN_347; // @[loaf.scala 176:26]
  wire  _GEN_352; // @[loaf.scala 176:26]
  wire  _GEN_357; // @[loaf.scala 176:26]
  wire  _GEN_362; // @[loaf.scala 176:26]
  wire  _GEN_367; // @[loaf.scala 176:26]
  wire  _GEN_372; // @[loaf.scala 176:26]
  wire  _GEN_377; // @[loaf.scala 176:26]
  wire  _GEN_382; // @[loaf.scala 176:26]
  wire  _GEN_387; // @[loaf.scala 176:26]
  wire  _GEN_392; // @[loaf.scala 176:26]
  wire  _GEN_397; // @[loaf.scala 176:26]
  wire  _GEN_402; // @[loaf.scala 176:26]
  wire  _GEN_407; // @[loaf.scala 176:26]
  wire  _GEN_412; // @[loaf.scala 176:26]
  wire  _GEN_417; // @[loaf.scala 176:26]
  wire  _GEN_422; // @[loaf.scala 176:26]
  wire  _GEN_427; // @[loaf.scala 176:26]
  wire  _GEN_432; // @[loaf.scala 176:26]
  wire  _GEN_437; // @[loaf.scala 176:26]
  wire  _GEN_442; // @[loaf.scala 176:26]
  wire  _GEN_447; // @[loaf.scala 176:26]
  wire  _GEN_452; // @[loaf.scala 176:26]
  wire  _GEN_457; // @[loaf.scala 176:26]
  wire  _GEN_462; // @[loaf.scala 176:26]
  wire  _GEN_467; // @[loaf.scala 176:26]
  wire  _GEN_472; // @[loaf.scala 176:26]
  wire  _GEN_477; // @[loaf.scala 176:26]
  wire  _GEN_482; // @[loaf.scala 176:26]
  wire  _GEN_487; // @[loaf.scala 176:26]
  wire  _GEN_492; // @[loaf.scala 176:26]
  wire  _GEN_497; // @[loaf.scala 176:26]
  wire  _GEN_502; // @[loaf.scala 176:26]
  wire  _GEN_507; // @[loaf.scala 176:26]
  wire  _GEN_512; // @[loaf.scala 176:26]
  wire  _GEN_517; // @[loaf.scala 176:26]
  wire  _GEN_522; // @[loaf.scala 176:26]
  wire  _GEN_527; // @[loaf.scala 176:26]
  wire  _GEN_532; // @[loaf.scala 176:26]
  wire  _GEN_537; // @[loaf.scala 176:26]
  wire  _GEN_542; // @[loaf.scala 176:26]
  wire  _GEN_547; // @[loaf.scala 176:26]
  wire  _GEN_552; // @[loaf.scala 176:26]
  wire  _GEN_557; // @[loaf.scala 176:26]
  wire  _GEN_562; // @[loaf.scala 176:26]
  wire  _GEN_567; // @[loaf.scala 176:26]
  wire  _GEN_572; // @[loaf.scala 176:26]
  wire  _GEN_577; // @[loaf.scala 176:26]
  wire  _GEN_582; // @[loaf.scala 176:26]
  wire  _GEN_587; // @[loaf.scala 176:26]
  wire  _GEN_592; // @[loaf.scala 176:26]
  wire  _GEN_597; // @[loaf.scala 176:26]
  wire  _GEN_602; // @[loaf.scala 176:26]
  wire  _GEN_607; // @[loaf.scala 176:26]
  wire  _GEN_612; // @[loaf.scala 176:26]
  wire  _GEN_617; // @[loaf.scala 176:26]
  wire  _GEN_622; // @[loaf.scala 176:26]
  wire  _GEN_627; // @[loaf.scala 176:26]
  wire  _GEN_632; // @[loaf.scala 176:26]
  wire  _GEN_637; // @[loaf.scala 176:26]
  wire [2:0] _T_388; // @[loaf.scala 193:19]
  wire [1:0] _T_389; // @[loaf.scala 195:28]
  wire [2:0] _T_390; // @[loaf.scala 197:19]
  wire [1:0] _T_391; // @[loaf.scala 199:28]
  wire [4:0] _T_392; // @[loaf.scala 201:32]
  wire [3:0] _T_393; // @[loaf.scala 201:68]
  wire [4:0] _GEN_4793; // @[loaf.scala 201:59]
  wire [4:0] _T_395; // @[loaf.scala 201:59]
  wire [4:0] _GEN_4794; // @[loaf.scala 201:92]
  wire [4:0] _T_397; // @[loaf.scala 201:92]
  wire  _T_398; // @[loaf.scala 209:25]
  wire [4:0] _T_400; // @[loaf.scala 210:30]
  wire  _T_401; // @[loaf.scala 213:27]
  wire [4:0] _T_403; // @[loaf.scala 214:32]
  wire  _GEN_647; // @[loaf.scala 185:26]
  wire  _GEN_658; // @[loaf.scala 174:40]
  wire  _GEN_663; // @[loaf.scala 174:40]
  wire  _GEN_668; // @[loaf.scala 174:40]
  wire  _GEN_673; // @[loaf.scala 174:40]
  wire  _GEN_678; // @[loaf.scala 174:40]
  wire  _GEN_683; // @[loaf.scala 174:40]
  wire  _GEN_688; // @[loaf.scala 174:40]
  wire  _GEN_693; // @[loaf.scala 174:40]
  wire  _GEN_698; // @[loaf.scala 174:40]
  wire  _GEN_703; // @[loaf.scala 174:40]
  wire  _GEN_708; // @[loaf.scala 174:40]
  wire  _GEN_713; // @[loaf.scala 174:40]
  wire  _GEN_718; // @[loaf.scala 174:40]
  wire  _GEN_723; // @[loaf.scala 174:40]
  wire  _GEN_728; // @[loaf.scala 174:40]
  wire  _GEN_733; // @[loaf.scala 174:40]
  wire  _GEN_738; // @[loaf.scala 174:40]
  wire  _GEN_743; // @[loaf.scala 174:40]
  wire  _GEN_748; // @[loaf.scala 174:40]
  wire  _GEN_753; // @[loaf.scala 174:40]
  wire  _GEN_758; // @[loaf.scala 174:40]
  wire  _GEN_763; // @[loaf.scala 174:40]
  wire  _GEN_768; // @[loaf.scala 174:40]
  wire  _GEN_773; // @[loaf.scala 174:40]
  wire  _GEN_778; // @[loaf.scala 174:40]
  wire  _GEN_783; // @[loaf.scala 174:40]
  wire  _GEN_788; // @[loaf.scala 174:40]
  wire  _GEN_793; // @[loaf.scala 174:40]
  wire  _GEN_798; // @[loaf.scala 174:40]
  wire  _GEN_803; // @[loaf.scala 174:40]
  wire  _GEN_808; // @[loaf.scala 174:40]
  wire  _GEN_813; // @[loaf.scala 174:40]
  wire  _GEN_818; // @[loaf.scala 174:40]
  wire  _GEN_823; // @[loaf.scala 174:40]
  wire  _GEN_828; // @[loaf.scala 174:40]
  wire  _GEN_833; // @[loaf.scala 174:40]
  wire  _GEN_838; // @[loaf.scala 174:40]
  wire  _GEN_843; // @[loaf.scala 174:40]
  wire  _GEN_848; // @[loaf.scala 174:40]
  wire  _GEN_853; // @[loaf.scala 174:40]
  wire  _GEN_858; // @[loaf.scala 174:40]
  wire  _GEN_863; // @[loaf.scala 174:40]
  wire  _GEN_868; // @[loaf.scala 174:40]
  wire  _GEN_873; // @[loaf.scala 174:40]
  wire  _GEN_878; // @[loaf.scala 174:40]
  wire  _GEN_883; // @[loaf.scala 174:40]
  wire  _GEN_888; // @[loaf.scala 174:40]
  wire  _GEN_893; // @[loaf.scala 174:40]
  wire  _GEN_898; // @[loaf.scala 174:40]
  wire  _GEN_903; // @[loaf.scala 174:40]
  wire  _GEN_908; // @[loaf.scala 174:40]
  wire  _GEN_913; // @[loaf.scala 174:40]
  wire  _GEN_918; // @[loaf.scala 174:40]
  wire  _GEN_923; // @[loaf.scala 174:40]
  wire  _GEN_928; // @[loaf.scala 174:40]
  wire  _GEN_933; // @[loaf.scala 174:40]
  wire  _GEN_938; // @[loaf.scala 174:40]
  wire  _GEN_943; // @[loaf.scala 174:40]
  wire  _GEN_948; // @[loaf.scala 174:40]
  wire  _GEN_953; // @[loaf.scala 174:40]
  wire  _GEN_958; // @[loaf.scala 174:40]
  wire  _GEN_963; // @[loaf.scala 174:40]
  wire  _GEN_968; // @[loaf.scala 174:40]
  wire  _GEN_973; // @[loaf.scala 174:40]
  wire  _GEN_978; // @[loaf.scala 174:40]
  wire  _GEN_989; // @[loaf.scala 172:25]
  wire  _GEN_994; // @[loaf.scala 172:25]
  wire  _GEN_999; // @[loaf.scala 172:25]
  wire  _GEN_1004; // @[loaf.scala 172:25]
  wire  _GEN_1009; // @[loaf.scala 172:25]
  wire  _GEN_1014; // @[loaf.scala 172:25]
  wire  _GEN_1019; // @[loaf.scala 172:25]
  wire  _GEN_1024; // @[loaf.scala 172:25]
  wire  _GEN_1029; // @[loaf.scala 172:25]
  wire  _GEN_1034; // @[loaf.scala 172:25]
  wire  _GEN_1039; // @[loaf.scala 172:25]
  wire  _GEN_1044; // @[loaf.scala 172:25]
  wire  _GEN_1049; // @[loaf.scala 172:25]
  wire  _GEN_1054; // @[loaf.scala 172:25]
  wire  _GEN_1059; // @[loaf.scala 172:25]
  wire  _GEN_1064; // @[loaf.scala 172:25]
  wire  _GEN_1069; // @[loaf.scala 172:25]
  wire  _GEN_1074; // @[loaf.scala 172:25]
  wire  _GEN_1079; // @[loaf.scala 172:25]
  wire  _GEN_1084; // @[loaf.scala 172:25]
  wire  _GEN_1089; // @[loaf.scala 172:25]
  wire  _GEN_1094; // @[loaf.scala 172:25]
  wire  _GEN_1099; // @[loaf.scala 172:25]
  wire  _GEN_1104; // @[loaf.scala 172:25]
  wire  _GEN_1109; // @[loaf.scala 172:25]
  wire  _GEN_1114; // @[loaf.scala 172:25]
  wire  _GEN_1119; // @[loaf.scala 172:25]
  wire  _GEN_1124; // @[loaf.scala 172:25]
  wire  _GEN_1129; // @[loaf.scala 172:25]
  wire  _GEN_1134; // @[loaf.scala 172:25]
  wire  _GEN_1139; // @[loaf.scala 172:25]
  wire  _GEN_1144; // @[loaf.scala 172:25]
  wire  _GEN_1149; // @[loaf.scala 172:25]
  wire  _GEN_1154; // @[loaf.scala 172:25]
  wire  _GEN_1159; // @[loaf.scala 172:25]
  wire  _GEN_1164; // @[loaf.scala 172:25]
  wire  _GEN_1169; // @[loaf.scala 172:25]
  wire  _GEN_1174; // @[loaf.scala 172:25]
  wire  _GEN_1179; // @[loaf.scala 172:25]
  wire  _GEN_1184; // @[loaf.scala 172:25]
  wire  _GEN_1189; // @[loaf.scala 172:25]
  wire  _GEN_1194; // @[loaf.scala 172:25]
  wire  _GEN_1199; // @[loaf.scala 172:25]
  wire  _GEN_1204; // @[loaf.scala 172:25]
  wire  _GEN_1209; // @[loaf.scala 172:25]
  wire  _GEN_1214; // @[loaf.scala 172:25]
  wire  _GEN_1219; // @[loaf.scala 172:25]
  wire  _GEN_1224; // @[loaf.scala 172:25]
  wire  _GEN_1229; // @[loaf.scala 172:25]
  wire  _GEN_1234; // @[loaf.scala 172:25]
  wire  _GEN_1239; // @[loaf.scala 172:25]
  wire  _GEN_1244; // @[loaf.scala 172:25]
  wire  _GEN_1249; // @[loaf.scala 172:25]
  wire  _GEN_1254; // @[loaf.scala 172:25]
  wire  _GEN_1259; // @[loaf.scala 172:25]
  wire  _GEN_1264; // @[loaf.scala 172:25]
  wire  _GEN_1269; // @[loaf.scala 172:25]
  wire  _GEN_1274; // @[loaf.scala 172:25]
  wire  _GEN_1279; // @[loaf.scala 172:25]
  wire  _GEN_1284; // @[loaf.scala 172:25]
  wire  _GEN_1289; // @[loaf.scala 172:25]
  wire  _GEN_1294; // @[loaf.scala 172:25]
  wire  _GEN_1299; // @[loaf.scala 172:25]
  wire  _GEN_1304; // @[loaf.scala 172:25]
  wire  _GEN_1309; // @[loaf.scala 172:25]
  reg  _T_405; // @[tsr.scala 8:42]
  reg [31:0] _RAND_473;
  reg  _T_406; // @[tsr.scala 8:42]
  reg [31:0] _RAND_474;
  reg  _T_407; // @[tsr.scala 8:42]
  reg [31:0] _RAND_475;
  reg  _T_408; // @[tsr.scala 8:42]
  reg [31:0] _RAND_476;
  reg  _T_409; // @[tsr.scala 8:42]
  reg [31:0] _RAND_477;
  reg  _T_410; // @[tsr.scala 8:42]
  reg [31:0] _RAND_478;
  reg  _T_411; // @[tsr.scala 8:42]
  reg [31:0] _RAND_479;
  reg  _T_412; // @[tsr.scala 8:42]
  reg [31:0] _RAND_480;
  reg  _T_413; // @[tsr.scala 8:42]
  reg [31:0] _RAND_481;
  reg  _T_414; // @[tsr.scala 8:42]
  reg [31:0] _RAND_482;
  reg  _T_415; // @[tsr.scala 8:42]
  reg [31:0] _RAND_483;
  reg  _T_416; // @[tsr.scala 8:42]
  reg [31:0] _RAND_484;
  reg  _T_417; // @[tsr.scala 8:42]
  reg [31:0] _RAND_485;
  reg  _T_418; // @[tsr.scala 8:42]
  reg [31:0] _RAND_486;
  reg  _T_421; // @[tsr.scala 8:42]
  reg [31:0] _RAND_487;
  reg  _T_422; // @[tsr.scala 8:42]
  reg [31:0] _RAND_488;
  reg  _T_423; // @[tsr.scala 8:42]
  reg [31:0] _RAND_489;
  reg  _T_424; // @[tsr.scala 8:42]
  reg [31:0] _RAND_490;
  reg  _T_425; // @[tsr.scala 8:42]
  reg [31:0] _RAND_491;
  reg  _T_426; // @[tsr.scala 8:42]
  reg [31:0] _RAND_492;
  reg  _T_427; // @[tsr.scala 8:42]
  reg [31:0] _RAND_493;
  reg  _T_428; // @[tsr.scala 8:42]
  reg [31:0] _RAND_494;
  reg  _T_429; // @[tsr.scala 8:42]
  reg [31:0] _RAND_495;
  reg  _T_430; // @[tsr.scala 8:42]
  reg [31:0] _RAND_496;
  reg  _T_431; // @[tsr.scala 8:42]
  reg [31:0] _RAND_497;
  reg  _T_432; // @[tsr.scala 8:42]
  reg [31:0] _RAND_498;
  reg  _T_433; // @[tsr.scala 8:42]
  reg [31:0] _RAND_499;
  reg  _T_434; // @[tsr.scala 8:42]
  reg [31:0] _RAND_500;
  reg  _T_437; // @[tsr.scala 8:42]
  reg [31:0] _RAND_501;
  reg  _T_438; // @[tsr.scala 8:42]
  reg [31:0] _RAND_502;
  reg  _T_439; // @[tsr.scala 8:42]
  reg [31:0] _RAND_503;
  reg  _T_440; // @[tsr.scala 8:42]
  reg [31:0] _RAND_504;
  reg  _T_441; // @[tsr.scala 8:42]
  reg [31:0] _RAND_505;
  reg  _T_442; // @[tsr.scala 8:42]
  reg [31:0] _RAND_506;
  reg  _T_443; // @[tsr.scala 8:42]
  reg [31:0] _RAND_507;
  reg  _T_444; // @[tsr.scala 8:42]
  reg [31:0] _RAND_508;
  reg  _T_445; // @[tsr.scala 8:42]
  reg [31:0] _RAND_509;
  reg  _T_446; // @[tsr.scala 8:42]
  reg [31:0] _RAND_510;
  reg  _T_447; // @[tsr.scala 8:42]
  reg [31:0] _RAND_511;
  reg  _T_448; // @[tsr.scala 8:42]
  reg [31:0] _RAND_512;
  wire  _T_450; // @[loaf.scala 234:22]
  wire  _T_451; // @[loaf.scala 234:19]
  wire  _T_452; // @[loaf.scala 236:24]
  wire  _T_453; // @[loaf.scala 244:34]
  wire  _T_454; // @[loaf.scala 244:47]
  wire  _T_455; // @[loaf.scala 244:42]
  wire  _T_456; // @[loaf.scala 244:59]
  wire  _T_457; // @[loaf.scala 244:79]
  wire  _T_458; // @[loaf.scala 244:90]
  wire  _T_459; // @[loaf.scala 244:87]
  wire  _T_460; // @[loaf.scala 244:73]
  wire  _T_461; // @[loaf.scala 244:55]
  wire  _T_462; // @[loaf.scala 246:14]
  wire  _T_463; // @[loaf.scala 246:32]
  wire  _T_465; // @[loaf.scala 248:46]
  wire  _T_466; // @[loaf.scala 248:43]
  wire  _T_468; // @[loaf.scala 249:47]
  wire  _T_469; // @[loaf.scala 249:42]
  wire  _T_471; // @[loaf.scala 249:61]
  wire  _T_474; // @[loaf.scala 250:43]
  wire  _T_476; // @[loaf.scala 250:56]
  wire  _GEN_1763; // @[loaf.scala 257:50]
  wire  _T_485; // @[loaf.scala 267:43]
  wire  _T_487; // @[loaf.scala 267:56]
  wire [4:0] _T_491; // @[loaf.scala 275:39]
  wire [3:0] _T_492; // @[loaf.scala 275:72]
  wire [4:0] _GEN_4795; // @[loaf.scala 275:66]
  wire [4:0] _T_494; // @[loaf.scala 275:66]
  wire [4:0] _GEN_4796; // @[loaf.scala 275:96]
  wire [31:0] _T_499;
  wire [15:0] _T_500; // @[loaf.scala 276:58]
  wire [15:0] _T_501; // @[loaf.scala 276:58]
  wire [31:0] _T_510;
  wire [15:0] _T_511; // @[loaf.scala 276:58]
  wire [15:0] _T_512; // @[loaf.scala 276:58]
  wire [31:0] _T_521;
  wire [15:0] _T_522; // @[loaf.scala 276:58]
  wire [15:0] _T_523; // @[loaf.scala 276:58]
  wire [31:0] _T_532;
  wire [15:0] _T_533; // @[loaf.scala 276:58]
  wire [15:0] _T_534; // @[loaf.scala 276:58]
  wire [31:0] _T_543;
  wire [15:0] _T_544; // @[loaf.scala 276:58]
  wire [15:0] _T_545; // @[loaf.scala 276:58]
  wire [31:0] _T_554;
  wire [15:0] _T_555; // @[loaf.scala 276:58]
  wire [15:0] _T_556; // @[loaf.scala 276:58]
  wire [31:0] _T_565;
  wire [15:0] _T_566; // @[loaf.scala 276:58]
  wire [15:0] _T_567; // @[loaf.scala 276:58]
  wire [31:0] _T_576;
  wire [15:0] _T_577; // @[loaf.scala 276:58]
  wire [15:0] _T_578; // @[loaf.scala 276:58]
  wire [31:0] _T_587;
  wire [15:0] _T_588; // @[loaf.scala 276:58]
  wire [15:0] _T_589; // @[loaf.scala 276:58]
  wire [31:0] _T_598;
  wire [15:0] _T_599; // @[loaf.scala 276:58]
  wire [15:0] _T_600; // @[loaf.scala 276:58]
  wire [31:0] _T_609;
  wire [15:0] _T_610; // @[loaf.scala 276:58]
  wire [15:0] _T_611; // @[loaf.scala 276:58]
  wire [31:0] _T_620;
  wire [15:0] _T_621; // @[loaf.scala 276:58]
  wire [15:0] _T_622; // @[loaf.scala 276:58]
  wire [31:0] _T_631;
  wire [15:0] _T_632; // @[loaf.scala 276:58]
  wire [15:0] _T_633; // @[loaf.scala 276:58]
  wire [31:0] _T_642;
  wire [15:0] _T_643; // @[loaf.scala 276:58]
  wire [15:0] _T_644; // @[loaf.scala 276:58]
  wire [31:0] _T_653;
  wire [15:0] _T_654; // @[loaf.scala 276:58]
  wire [15:0] _T_655; // @[loaf.scala 276:58]
  wire [31:0] _T_664;
  wire [15:0] _T_665; // @[loaf.scala 276:58]
  wire [15:0] _T_666; // @[loaf.scala 276:58]
  wire [31:0] _T_675;
  wire [15:0] _T_676; // @[loaf.scala 276:58]
  wire [15:0] _T_677; // @[loaf.scala 276:58]
  wire [31:0] _T_686;
  wire [15:0] _T_687; // @[loaf.scala 276:58]
  wire [15:0] _T_688; // @[loaf.scala 276:58]
  wire [31:0] _T_697;
  wire [15:0] _T_698; // @[loaf.scala 276:58]
  wire [15:0] _T_699; // @[loaf.scala 276:58]
  wire [31:0] _T_708;
  wire [15:0] _T_709; // @[loaf.scala 276:58]
  wire [15:0] _T_710; // @[loaf.scala 276:58]
  wire [31:0] _T_719;
  wire [15:0] _T_720; // @[loaf.scala 276:58]
  wire [15:0] _T_721; // @[loaf.scala 276:58]
  wire [31:0] _T_730;
  wire [15:0] _T_731; // @[loaf.scala 276:58]
  wire [15:0] _T_732; // @[loaf.scala 276:58]
  wire [31:0] _T_741;
  wire [15:0] _T_742; // @[loaf.scala 276:58]
  wire [15:0] _T_743; // @[loaf.scala 276:58]
  wire [31:0] _T_752;
  wire [15:0] _T_753; // @[loaf.scala 276:58]
  wire [15:0] _T_754; // @[loaf.scala 276:58]
  wire [31:0] _T_763;
  wire [15:0] _T_764; // @[loaf.scala 276:58]
  wire [15:0] _T_765; // @[loaf.scala 276:58]
  wire [31:0] _T_774;
  wire [15:0] _T_775; // @[loaf.scala 276:58]
  wire [15:0] _T_776; // @[loaf.scala 276:58]
  wire [31:0] _T_785;
  wire [15:0] _T_786; // @[loaf.scala 276:58]
  wire [15:0] _T_787; // @[loaf.scala 276:58]
  wire [31:0] _T_796;
  wire [15:0] _T_797; // @[loaf.scala 276:58]
  wire [15:0] _T_798; // @[loaf.scala 276:58]
  wire [31:0] _T_807;
  wire [15:0] _T_808; // @[loaf.scala 276:58]
  wire [15:0] _T_809; // @[loaf.scala 276:58]
  wire [31:0] _T_818;
  wire [15:0] _T_819; // @[loaf.scala 276:58]
  wire [15:0] _T_820; // @[loaf.scala 276:58]
  wire [31:0] _T_829;
  wire [15:0] _T_830; // @[loaf.scala 276:58]
  wire [15:0] _T_831; // @[loaf.scala 276:58]
  wire [31:0] _T_840;
  wire [15:0] _T_841; // @[loaf.scala 276:58]
  wire [15:0] _T_842; // @[loaf.scala 276:58]
  wire [31:0] _T_851;
  wire [15:0] _T_852; // @[loaf.scala 276:58]
  wire [15:0] _T_853; // @[loaf.scala 276:58]
  wire [31:0] _T_862;
  wire [15:0] _T_863; // @[loaf.scala 276:58]
  wire [15:0] _T_864; // @[loaf.scala 276:58]
  wire [31:0] _T_873;
  wire [15:0] _T_874; // @[loaf.scala 276:58]
  wire [15:0] _T_875; // @[loaf.scala 276:58]
  wire [31:0] _T_884;
  wire [15:0] _T_885; // @[loaf.scala 276:58]
  wire [15:0] _T_886; // @[loaf.scala 276:58]
  wire [31:0] _T_895;
  wire [15:0] _T_896; // @[loaf.scala 276:58]
  wire [15:0] _T_897; // @[loaf.scala 276:58]
  wire [31:0] _T_906;
  wire [15:0] _T_907; // @[loaf.scala 276:58]
  wire [15:0] _T_908; // @[loaf.scala 276:58]
  wire [31:0] _T_917;
  wire [15:0] _T_918; // @[loaf.scala 276:58]
  wire [15:0] _T_919; // @[loaf.scala 276:58]
  wire [31:0] _T_928;
  wire [15:0] _T_929; // @[loaf.scala 276:58]
  wire [15:0] _T_930; // @[loaf.scala 276:58]
  wire [31:0] _T_939;
  wire [15:0] _T_940; // @[loaf.scala 276:58]
  wire [15:0] _T_941; // @[loaf.scala 276:58]
  wire [31:0] _T_950;
  wire [15:0] _T_951; // @[loaf.scala 276:58]
  wire [15:0] _T_952; // @[loaf.scala 276:58]
  wire [31:0] _T_961;
  wire [15:0] _T_962; // @[loaf.scala 276:58]
  wire [15:0] _T_963; // @[loaf.scala 276:58]
  wire [31:0] _T_972;
  wire [15:0] _T_973; // @[loaf.scala 276:58]
  wire [15:0] _T_974; // @[loaf.scala 276:58]
  wire [31:0] _T_983;
  wire [15:0] _T_984; // @[loaf.scala 276:58]
  wire [15:0] _T_985; // @[loaf.scala 276:58]
  wire [31:0] _T_994;
  wire [15:0] _T_995; // @[loaf.scala 276:58]
  wire [15:0] _T_996; // @[loaf.scala 276:58]
  wire [31:0] _T_1005;
  wire [15:0] _T_1006; // @[loaf.scala 276:58]
  wire [15:0] _T_1007; // @[loaf.scala 276:58]
  wire [31:0] _T_1016;
  wire [15:0] _T_1017; // @[loaf.scala 276:58]
  wire [15:0] _T_1018; // @[loaf.scala 276:58]
  wire [31:0] _T_1027;
  wire [15:0] _T_1028; // @[loaf.scala 276:58]
  wire [15:0] _T_1029; // @[loaf.scala 276:58]
  wire [31:0] _T_1038;
  wire [15:0] _T_1039; // @[loaf.scala 276:58]
  wire [15:0] _T_1040; // @[loaf.scala 276:58]
  wire [31:0] _T_1049;
  wire [15:0] _T_1050; // @[loaf.scala 276:58]
  wire [15:0] _T_1051; // @[loaf.scala 276:58]
  wire [31:0] _T_1060;
  wire [15:0] _T_1061; // @[loaf.scala 276:58]
  wire [15:0] _T_1062; // @[loaf.scala 276:58]
  wire [31:0] _T_1071;
  wire [15:0] _T_1072; // @[loaf.scala 276:58]
  wire [15:0] _T_1073; // @[loaf.scala 276:58]
  wire [31:0] _T_1082;
  wire [15:0] _T_1083; // @[loaf.scala 276:58]
  wire [15:0] _T_1084; // @[loaf.scala 276:58]
  wire [31:0] _T_1093;
  wire [15:0] _T_1094; // @[loaf.scala 276:58]
  wire [15:0] _T_1095; // @[loaf.scala 276:58]
  wire [31:0] _T_1104;
  wire [15:0] _T_1105; // @[loaf.scala 276:58]
  wire [15:0] _T_1106; // @[loaf.scala 276:58]
  wire [31:0] _T_1115;
  wire [15:0] _T_1116; // @[loaf.scala 276:58]
  wire [15:0] _T_1117; // @[loaf.scala 276:58]
  wire [31:0] _T_1126;
  wire [15:0] _T_1127; // @[loaf.scala 276:58]
  wire [15:0] _T_1128; // @[loaf.scala 276:58]
  wire [31:0] _T_1137;
  wire [15:0] _T_1138; // @[loaf.scala 276:58]
  wire [15:0] _T_1139; // @[loaf.scala 276:58]
  wire [31:0] _T_1148;
  wire [15:0] _T_1149; // @[loaf.scala 276:58]
  wire [15:0] _T_1150; // @[loaf.scala 276:58]
  wire [31:0] _T_1159;
  wire [15:0] _T_1160; // @[loaf.scala 276:58]
  wire [15:0] _T_1161; // @[loaf.scala 276:58]
  wire [31:0] _T_1170;
  wire [15:0] _T_1171; // @[loaf.scala 276:58]
  wire [15:0] _T_1172; // @[loaf.scala 276:58]
  wire [31:0] _T_1181;
  wire [15:0] _T_1182; // @[loaf.scala 276:58]
  wire [15:0] _T_1183; // @[loaf.scala 276:58]
  wire [31:0] _T_1192;
  wire [15:0] _T_1193; // @[loaf.scala 276:58]
  wire [15:0] _T_1194; // @[loaf.scala 276:58]
  wire  _T_1196; // @[loaf.scala 292:22]
  wire [15:0] _T_1198; // @[loaf.scala 294:33]
  wire  _T_1200; // @[loaf.scala 295:21]
  wire [15:0] _T_1202; // @[loaf.scala 295:34]
  wire  _T_1204; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2003; // @[loaf.scala 298:37]
  wire [25:0] _T_1205; // @[loaf.scala 302:38]
  wire [21:0] _T_1206; // @[loaf.scala 316:29]
  wire  _T_1208; // @[loaf.scala 292:22]
  wire [15:0] _T_1210; // @[loaf.scala 294:33]
  wire  _T_1212; // @[loaf.scala 295:21]
  wire [15:0] _T_1214; // @[loaf.scala 295:34]
  wire  _T_1216; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2006; // @[loaf.scala 298:37]
  wire [25:0] _T_1217; // @[loaf.scala 302:38]
  wire [21:0] _T_1218; // @[loaf.scala 316:29]
  wire  _T_1220; // @[loaf.scala 292:22]
  wire [15:0] _T_1222; // @[loaf.scala 294:33]
  wire  _T_1224; // @[loaf.scala 295:21]
  wire [15:0] _T_1226; // @[loaf.scala 295:34]
  wire  _T_1228; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2009; // @[loaf.scala 298:37]
  wire [25:0] _T_1229; // @[loaf.scala 302:38]
  wire [21:0] _T_1230; // @[loaf.scala 316:29]
  wire  _T_1232; // @[loaf.scala 292:22]
  wire [15:0] _T_1234; // @[loaf.scala 294:33]
  wire  _T_1236; // @[loaf.scala 295:21]
  wire [15:0] _T_1238; // @[loaf.scala 295:34]
  wire  _T_1240; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2012; // @[loaf.scala 298:37]
  wire [25:0] _T_1241; // @[loaf.scala 302:38]
  wire [21:0] _T_1242; // @[loaf.scala 316:29]
  wire  _T_1244; // @[loaf.scala 292:22]
  wire [15:0] _T_1246; // @[loaf.scala 294:33]
  wire  _T_1248; // @[loaf.scala 295:21]
  wire [15:0] _T_1250; // @[loaf.scala 295:34]
  wire  _T_1252; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2015; // @[loaf.scala 298:37]
  wire [25:0] _T_1253; // @[loaf.scala 302:38]
  wire [21:0] _T_1254; // @[loaf.scala 316:29]
  wire  _T_1256; // @[loaf.scala 292:22]
  wire [15:0] _T_1258; // @[loaf.scala 294:33]
  wire  _T_1260; // @[loaf.scala 295:21]
  wire [15:0] _T_1262; // @[loaf.scala 295:34]
  wire  _T_1264; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2018; // @[loaf.scala 298:37]
  wire [25:0] _T_1265; // @[loaf.scala 302:38]
  wire [21:0] _T_1266; // @[loaf.scala 316:29]
  wire  _T_1268; // @[loaf.scala 292:22]
  wire [15:0] _T_1270; // @[loaf.scala 294:33]
  wire  _T_1272; // @[loaf.scala 295:21]
  wire [15:0] _T_1274; // @[loaf.scala 295:34]
  wire  _T_1276; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2021; // @[loaf.scala 298:37]
  wire [25:0] _T_1277; // @[loaf.scala 302:38]
  wire [21:0] _T_1278; // @[loaf.scala 316:29]
  wire  _T_1280; // @[loaf.scala 292:22]
  wire [15:0] _T_1282; // @[loaf.scala 294:33]
  wire  _T_1284; // @[loaf.scala 295:21]
  wire [15:0] _T_1286; // @[loaf.scala 295:34]
  wire  _T_1288; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2024; // @[loaf.scala 298:37]
  wire [25:0] _T_1289; // @[loaf.scala 302:38]
  wire [21:0] _T_1290; // @[loaf.scala 316:29]
  wire  _T_1292; // @[loaf.scala 327:24]
  wire [21:0] _GEN_2025; // @[loaf.scala 327:29]
  wire  _T_1294; // @[loaf.scala 327:24]
  wire [21:0] _GEN_2026; // @[loaf.scala 327:29]
  wire  _T_1296; // @[loaf.scala 327:24]
  wire [21:0] _GEN_2027; // @[loaf.scala 327:29]
  wire  _T_1298; // @[loaf.scala 327:24]
  wire [21:0] _GEN_2028; // @[loaf.scala 327:29]
  wire  _T_1300; // @[loaf.scala 327:24]
  wire  _T_1302; // @[loaf.scala 327:24]
  wire  _T_1304; // @[loaf.scala 327:24]
  wire  _T_1306; // @[loaf.scala 354:43]
  wire  _T_1307; // @[loaf.scala 354:35]
  wire  _T_1309; // @[loaf.scala 292:22]
  wire [15:0] _T_1311; // @[loaf.scala 294:33]
  wire  _T_1313; // @[loaf.scala 295:21]
  wire [15:0] _T_1315; // @[loaf.scala 295:34]
  wire  _T_1317; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2035; // @[loaf.scala 298:37]
  wire [21:0] _T_1319; // @[loaf.scala 316:29]
  wire  _T_1321; // @[loaf.scala 292:22]
  wire [15:0] _T_1323; // @[loaf.scala 294:33]
  wire  _T_1325; // @[loaf.scala 295:21]
  wire [15:0] _T_1327; // @[loaf.scala 295:34]
  wire  _T_1329; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2038; // @[loaf.scala 298:37]
  wire [21:0] _T_1331; // @[loaf.scala 316:29]
  wire  _T_1333; // @[loaf.scala 292:22]
  wire [15:0] _T_1335; // @[loaf.scala 294:33]
  wire  _T_1337; // @[loaf.scala 295:21]
  wire [15:0] _T_1339; // @[loaf.scala 295:34]
  wire  _T_1341; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2041; // @[loaf.scala 298:37]
  wire [21:0] _T_1343; // @[loaf.scala 316:29]
  wire  _T_1345; // @[loaf.scala 292:22]
  wire [15:0] _T_1347; // @[loaf.scala 294:33]
  wire  _T_1349; // @[loaf.scala 295:21]
  wire [15:0] _T_1351; // @[loaf.scala 295:34]
  wire  _T_1353; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2044; // @[loaf.scala 298:37]
  wire [21:0] _T_1355; // @[loaf.scala 316:29]
  wire  _T_1357; // @[loaf.scala 292:22]
  wire [15:0] _T_1359; // @[loaf.scala 294:33]
  wire  _T_1361; // @[loaf.scala 295:21]
  wire [15:0] _T_1363; // @[loaf.scala 295:34]
  wire  _T_1365; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2047; // @[loaf.scala 298:37]
  wire [21:0] _T_1367; // @[loaf.scala 316:29]
  wire  _T_1369; // @[loaf.scala 292:22]
  wire [15:0] _T_1371; // @[loaf.scala 294:33]
  wire  _T_1373; // @[loaf.scala 295:21]
  wire [15:0] _T_1375; // @[loaf.scala 295:34]
  wire  _T_1377; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2050; // @[loaf.scala 298:37]
  wire [21:0] _T_1379; // @[loaf.scala 316:29]
  wire  _T_1381; // @[loaf.scala 292:22]
  wire [15:0] _T_1383; // @[loaf.scala 294:33]
  wire  _T_1385; // @[loaf.scala 295:21]
  wire [15:0] _T_1387; // @[loaf.scala 295:34]
  wire  _T_1389; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2053; // @[loaf.scala 298:37]
  wire [21:0] _T_1391; // @[loaf.scala 316:29]
  wire  _T_1393; // @[loaf.scala 292:22]
  wire [15:0] _T_1395; // @[loaf.scala 294:33]
  wire  _T_1397; // @[loaf.scala 295:21]
  wire [15:0] _T_1399; // @[loaf.scala 295:34]
  wire  _T_1401; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2056; // @[loaf.scala 298:37]
  wire [21:0] _T_1403; // @[loaf.scala 316:29]
  wire  _T_1405; // @[loaf.scala 327:24]
  wire [21:0] _GEN_2057; // @[loaf.scala 327:29]
  wire  _T_1407; // @[loaf.scala 327:24]
  wire [21:0] _GEN_2058; // @[loaf.scala 327:29]
  wire  _T_1409; // @[loaf.scala 327:24]
  wire [21:0] _GEN_2059; // @[loaf.scala 327:29]
  wire  _T_1411; // @[loaf.scala 327:24]
  wire [21:0] _GEN_2060; // @[loaf.scala 327:29]
  wire  _T_1413; // @[loaf.scala 327:24]
  wire  _T_1415; // @[loaf.scala 327:24]
  wire  _T_1417; // @[loaf.scala 327:24]
  wire  _T_1419; // @[loaf.scala 354:43]
  wire  _T_1420; // @[loaf.scala 354:35]
  wire  _T_1422; // @[loaf.scala 292:22]
  wire [15:0] _T_1424; // @[loaf.scala 294:33]
  wire  _T_1426; // @[loaf.scala 295:21]
  wire [15:0] _T_1428; // @[loaf.scala 295:34]
  wire  _T_1430; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2067; // @[loaf.scala 298:37]
  wire [21:0] _T_1432; // @[loaf.scala 316:29]
  wire  _T_1434; // @[loaf.scala 292:22]
  wire [15:0] _T_1436; // @[loaf.scala 294:33]
  wire  _T_1438; // @[loaf.scala 295:21]
  wire [15:0] _T_1440; // @[loaf.scala 295:34]
  wire  _T_1442; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2070; // @[loaf.scala 298:37]
  wire [21:0] _T_1444; // @[loaf.scala 316:29]
  wire  _T_1446; // @[loaf.scala 292:22]
  wire [15:0] _T_1448; // @[loaf.scala 294:33]
  wire  _T_1450; // @[loaf.scala 295:21]
  wire [15:0] _T_1452; // @[loaf.scala 295:34]
  wire  _T_1454; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2073; // @[loaf.scala 298:37]
  wire [21:0] _T_1456; // @[loaf.scala 316:29]
  wire  _T_1458; // @[loaf.scala 292:22]
  wire [15:0] _T_1460; // @[loaf.scala 294:33]
  wire  _T_1462; // @[loaf.scala 295:21]
  wire [15:0] _T_1464; // @[loaf.scala 295:34]
  wire  _T_1466; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2076; // @[loaf.scala 298:37]
  wire [21:0] _T_1468; // @[loaf.scala 316:29]
  wire  _T_1470; // @[loaf.scala 292:22]
  wire [15:0] _T_1472; // @[loaf.scala 294:33]
  wire  _T_1474; // @[loaf.scala 295:21]
  wire [15:0] _T_1476; // @[loaf.scala 295:34]
  wire  _T_1478; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2079; // @[loaf.scala 298:37]
  wire [21:0] _T_1480; // @[loaf.scala 316:29]
  wire  _T_1482; // @[loaf.scala 292:22]
  wire [15:0] _T_1484; // @[loaf.scala 294:33]
  wire  _T_1486; // @[loaf.scala 295:21]
  wire [15:0] _T_1488; // @[loaf.scala 295:34]
  wire  _T_1490; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2082; // @[loaf.scala 298:37]
  wire [21:0] _T_1492; // @[loaf.scala 316:29]
  wire  _T_1494; // @[loaf.scala 292:22]
  wire [15:0] _T_1496; // @[loaf.scala 294:33]
  wire  _T_1498; // @[loaf.scala 295:21]
  wire [15:0] _T_1500; // @[loaf.scala 295:34]
  wire  _T_1502; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2085; // @[loaf.scala 298:37]
  wire [21:0] _T_1504; // @[loaf.scala 316:29]
  wire  _T_1506; // @[loaf.scala 292:22]
  wire [15:0] _T_1508; // @[loaf.scala 294:33]
  wire  _T_1510; // @[loaf.scala 295:21]
  wire [15:0] _T_1512; // @[loaf.scala 295:34]
  wire  _T_1514; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2088; // @[loaf.scala 298:37]
  wire [21:0] _T_1516; // @[loaf.scala 316:29]
  wire  _T_1518; // @[loaf.scala 327:24]
  wire [21:0] _GEN_2089; // @[loaf.scala 327:29]
  wire  _T_1520; // @[loaf.scala 327:24]
  wire [21:0] _GEN_2090; // @[loaf.scala 327:29]
  wire  _T_1522; // @[loaf.scala 327:24]
  wire [21:0] _GEN_2091; // @[loaf.scala 327:29]
  wire  _T_1524; // @[loaf.scala 327:24]
  wire [21:0] _GEN_2092; // @[loaf.scala 327:29]
  wire  _T_1526; // @[loaf.scala 327:24]
  wire  _T_1528; // @[loaf.scala 327:24]
  wire  _T_1530; // @[loaf.scala 327:24]
  wire  _T_1532; // @[loaf.scala 354:43]
  wire  _T_1533; // @[loaf.scala 354:35]
  wire  _T_1535; // @[loaf.scala 292:22]
  wire [15:0] _T_1537; // @[loaf.scala 294:33]
  wire  _T_1539; // @[loaf.scala 295:21]
  wire [15:0] _T_1541; // @[loaf.scala 295:34]
  wire  _T_1543; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2099; // @[loaf.scala 298:37]
  wire [21:0] _T_1545; // @[loaf.scala 316:29]
  wire  _T_1547; // @[loaf.scala 292:22]
  wire [15:0] _T_1549; // @[loaf.scala 294:33]
  wire  _T_1551; // @[loaf.scala 295:21]
  wire [15:0] _T_1553; // @[loaf.scala 295:34]
  wire  _T_1555; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2102; // @[loaf.scala 298:37]
  wire [21:0] _T_1557; // @[loaf.scala 316:29]
  wire  _T_1559; // @[loaf.scala 292:22]
  wire [15:0] _T_1561; // @[loaf.scala 294:33]
  wire  _T_1563; // @[loaf.scala 295:21]
  wire [15:0] _T_1565; // @[loaf.scala 295:34]
  wire  _T_1567; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2105; // @[loaf.scala 298:37]
  wire [21:0] _T_1569; // @[loaf.scala 316:29]
  wire  _T_1571; // @[loaf.scala 292:22]
  wire [15:0] _T_1573; // @[loaf.scala 294:33]
  wire  _T_1575; // @[loaf.scala 295:21]
  wire [15:0] _T_1577; // @[loaf.scala 295:34]
  wire  _T_1579; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2108; // @[loaf.scala 298:37]
  wire [21:0] _T_1581; // @[loaf.scala 316:29]
  wire  _T_1583; // @[loaf.scala 292:22]
  wire [15:0] _T_1585; // @[loaf.scala 294:33]
  wire  _T_1587; // @[loaf.scala 295:21]
  wire [15:0] _T_1589; // @[loaf.scala 295:34]
  wire  _T_1591; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2111; // @[loaf.scala 298:37]
  wire [21:0] _T_1593; // @[loaf.scala 316:29]
  wire  _T_1595; // @[loaf.scala 292:22]
  wire [15:0] _T_1597; // @[loaf.scala 294:33]
  wire  _T_1599; // @[loaf.scala 295:21]
  wire [15:0] _T_1601; // @[loaf.scala 295:34]
  wire  _T_1603; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2114; // @[loaf.scala 298:37]
  wire [21:0] _T_1605; // @[loaf.scala 316:29]
  wire  _T_1607; // @[loaf.scala 292:22]
  wire [15:0] _T_1609; // @[loaf.scala 294:33]
  wire  _T_1611; // @[loaf.scala 295:21]
  wire [15:0] _T_1613; // @[loaf.scala 295:34]
  wire  _T_1615; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2117; // @[loaf.scala 298:37]
  wire [21:0] _T_1617; // @[loaf.scala 316:29]
  wire  _T_1619; // @[loaf.scala 292:22]
  wire [15:0] _T_1621; // @[loaf.scala 294:33]
  wire  _T_1623; // @[loaf.scala 295:21]
  wire [15:0] _T_1625; // @[loaf.scala 295:34]
  wire  _T_1627; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2120; // @[loaf.scala 298:37]
  wire [21:0] _T_1629; // @[loaf.scala 316:29]
  wire  _T_1631; // @[loaf.scala 327:24]
  wire [21:0] _GEN_2121; // @[loaf.scala 327:29]
  wire  _T_1633; // @[loaf.scala 327:24]
  wire [21:0] _GEN_2122; // @[loaf.scala 327:29]
  wire  _T_1635; // @[loaf.scala 327:24]
  wire [21:0] _GEN_2123; // @[loaf.scala 327:29]
  wire  _T_1637; // @[loaf.scala 327:24]
  wire [21:0] _GEN_2124; // @[loaf.scala 327:29]
  wire  _T_1639; // @[loaf.scala 327:24]
  wire  _T_1641; // @[loaf.scala 327:24]
  wire  _T_1643; // @[loaf.scala 327:24]
  wire  _T_1645; // @[loaf.scala 354:43]
  wire  _T_1646; // @[loaf.scala 354:35]
  wire  _T_1648; // @[loaf.scala 292:22]
  wire [15:0] _T_1650; // @[loaf.scala 294:33]
  wire  _T_1652; // @[loaf.scala 295:21]
  wire [15:0] _T_1654; // @[loaf.scala 295:34]
  wire  _T_1656; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2131; // @[loaf.scala 298:37]
  wire [21:0] _T_1658; // @[loaf.scala 316:29]
  wire  _T_1660; // @[loaf.scala 292:22]
  wire [15:0] _T_1662; // @[loaf.scala 294:33]
  wire  _T_1664; // @[loaf.scala 295:21]
  wire [15:0] _T_1666; // @[loaf.scala 295:34]
  wire  _T_1668; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2134; // @[loaf.scala 298:37]
  wire [21:0] _T_1670; // @[loaf.scala 316:29]
  wire  _T_1672; // @[loaf.scala 292:22]
  wire [15:0] _T_1674; // @[loaf.scala 294:33]
  wire  _T_1676; // @[loaf.scala 295:21]
  wire [15:0] _T_1678; // @[loaf.scala 295:34]
  wire  _T_1680; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2137; // @[loaf.scala 298:37]
  wire [21:0] _T_1682; // @[loaf.scala 316:29]
  wire  _T_1684; // @[loaf.scala 292:22]
  wire [15:0] _T_1686; // @[loaf.scala 294:33]
  wire  _T_1688; // @[loaf.scala 295:21]
  wire [15:0] _T_1690; // @[loaf.scala 295:34]
  wire  _T_1692; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2140; // @[loaf.scala 298:37]
  wire [21:0] _T_1694; // @[loaf.scala 316:29]
  wire  _T_1696; // @[loaf.scala 292:22]
  wire [15:0] _T_1698; // @[loaf.scala 294:33]
  wire  _T_1700; // @[loaf.scala 295:21]
  wire [15:0] _T_1702; // @[loaf.scala 295:34]
  wire  _T_1704; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2143; // @[loaf.scala 298:37]
  wire [21:0] _T_1706; // @[loaf.scala 316:29]
  wire  _T_1708; // @[loaf.scala 292:22]
  wire [15:0] _T_1710; // @[loaf.scala 294:33]
  wire  _T_1712; // @[loaf.scala 295:21]
  wire [15:0] _T_1714; // @[loaf.scala 295:34]
  wire  _T_1716; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2146; // @[loaf.scala 298:37]
  wire [21:0] _T_1718; // @[loaf.scala 316:29]
  wire  _T_1720; // @[loaf.scala 292:22]
  wire [15:0] _T_1722; // @[loaf.scala 294:33]
  wire  _T_1724; // @[loaf.scala 295:21]
  wire [15:0] _T_1726; // @[loaf.scala 295:34]
  wire  _T_1728; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2149; // @[loaf.scala 298:37]
  wire [21:0] _T_1730; // @[loaf.scala 316:29]
  wire  _T_1732; // @[loaf.scala 292:22]
  wire [15:0] _T_1734; // @[loaf.scala 294:33]
  wire  _T_1736; // @[loaf.scala 295:21]
  wire [15:0] _T_1738; // @[loaf.scala 295:34]
  wire  _T_1740; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2152; // @[loaf.scala 298:37]
  wire [21:0] _T_1742; // @[loaf.scala 316:29]
  wire  _T_1744; // @[loaf.scala 327:24]
  wire [21:0] _GEN_2153; // @[loaf.scala 327:29]
  wire  _T_1746; // @[loaf.scala 327:24]
  wire [21:0] _GEN_2154; // @[loaf.scala 327:29]
  wire  _T_1748; // @[loaf.scala 327:24]
  wire [21:0] _GEN_2155; // @[loaf.scala 327:29]
  wire  _T_1750; // @[loaf.scala 327:24]
  wire [21:0] _GEN_2156; // @[loaf.scala 327:29]
  wire  _T_1752; // @[loaf.scala 327:24]
  wire  _T_1754; // @[loaf.scala 327:24]
  wire  _T_1756; // @[loaf.scala 327:24]
  wire  _T_1758; // @[loaf.scala 354:43]
  wire  _T_1759; // @[loaf.scala 354:35]
  wire  _T_1761; // @[loaf.scala 292:22]
  wire [15:0] _T_1763; // @[loaf.scala 294:33]
  wire  _T_1765; // @[loaf.scala 295:21]
  wire [15:0] _T_1767; // @[loaf.scala 295:34]
  wire  _T_1769; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2163; // @[loaf.scala 298:37]
  wire [21:0] _T_1771; // @[loaf.scala 316:29]
  wire  _T_1773; // @[loaf.scala 292:22]
  wire [15:0] _T_1775; // @[loaf.scala 294:33]
  wire  _T_1777; // @[loaf.scala 295:21]
  wire [15:0] _T_1779; // @[loaf.scala 295:34]
  wire  _T_1781; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2166; // @[loaf.scala 298:37]
  wire [21:0] _T_1783; // @[loaf.scala 316:29]
  wire  _T_1785; // @[loaf.scala 292:22]
  wire [15:0] _T_1787; // @[loaf.scala 294:33]
  wire  _T_1789; // @[loaf.scala 295:21]
  wire [15:0] _T_1791; // @[loaf.scala 295:34]
  wire  _T_1793; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2169; // @[loaf.scala 298:37]
  wire [21:0] _T_1795; // @[loaf.scala 316:29]
  wire  _T_1797; // @[loaf.scala 292:22]
  wire [15:0] _T_1799; // @[loaf.scala 294:33]
  wire  _T_1801; // @[loaf.scala 295:21]
  wire [15:0] _T_1803; // @[loaf.scala 295:34]
  wire  _T_1805; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2172; // @[loaf.scala 298:37]
  wire [21:0] _T_1807; // @[loaf.scala 316:29]
  wire  _T_1809; // @[loaf.scala 292:22]
  wire [15:0] _T_1811; // @[loaf.scala 294:33]
  wire  _T_1813; // @[loaf.scala 295:21]
  wire [15:0] _T_1815; // @[loaf.scala 295:34]
  wire  _T_1817; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2175; // @[loaf.scala 298:37]
  wire [21:0] _T_1819; // @[loaf.scala 316:29]
  wire  _T_1821; // @[loaf.scala 292:22]
  wire [15:0] _T_1823; // @[loaf.scala 294:33]
  wire  _T_1825; // @[loaf.scala 295:21]
  wire [15:0] _T_1827; // @[loaf.scala 295:34]
  wire  _T_1829; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2178; // @[loaf.scala 298:37]
  wire [21:0] _T_1831; // @[loaf.scala 316:29]
  wire  _T_1833; // @[loaf.scala 292:22]
  wire [15:0] _T_1835; // @[loaf.scala 294:33]
  wire  _T_1837; // @[loaf.scala 295:21]
  wire [15:0] _T_1839; // @[loaf.scala 295:34]
  wire  _T_1841; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2181; // @[loaf.scala 298:37]
  wire [21:0] _T_1843; // @[loaf.scala 316:29]
  wire  _T_1845; // @[loaf.scala 292:22]
  wire [15:0] _T_1847; // @[loaf.scala 294:33]
  wire  _T_1849; // @[loaf.scala 295:21]
  wire [15:0] _T_1851; // @[loaf.scala 295:34]
  wire  _T_1853; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2184; // @[loaf.scala 298:37]
  wire [21:0] _T_1855; // @[loaf.scala 316:29]
  wire  _T_1857; // @[loaf.scala 327:24]
  wire [21:0] _GEN_2185; // @[loaf.scala 327:29]
  wire  _T_1859; // @[loaf.scala 327:24]
  wire [21:0] _GEN_2186; // @[loaf.scala 327:29]
  wire  _T_1861; // @[loaf.scala 327:24]
  wire [21:0] _GEN_2187; // @[loaf.scala 327:29]
  wire  _T_1863; // @[loaf.scala 327:24]
  wire [21:0] _GEN_2188; // @[loaf.scala 327:29]
  wire  _T_1865; // @[loaf.scala 327:24]
  wire  _T_1867; // @[loaf.scala 327:24]
  wire  _T_1869; // @[loaf.scala 327:24]
  wire  _T_1871; // @[loaf.scala 354:43]
  wire  _T_1872; // @[loaf.scala 354:35]
  wire  _T_1874; // @[loaf.scala 292:22]
  wire [15:0] _T_1876; // @[loaf.scala 294:33]
  wire  _T_1878; // @[loaf.scala 295:21]
  wire [15:0] _T_1880; // @[loaf.scala 295:34]
  wire  _T_1882; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2195; // @[loaf.scala 298:37]
  wire [21:0] _T_1884; // @[loaf.scala 316:29]
  wire  _T_1886; // @[loaf.scala 292:22]
  wire [15:0] _T_1888; // @[loaf.scala 294:33]
  wire  _T_1890; // @[loaf.scala 295:21]
  wire [15:0] _T_1892; // @[loaf.scala 295:34]
  wire  _T_1894; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2198; // @[loaf.scala 298:37]
  wire [21:0] _T_1896; // @[loaf.scala 316:29]
  wire  _T_1898; // @[loaf.scala 292:22]
  wire [15:0] _T_1900; // @[loaf.scala 294:33]
  wire  _T_1902; // @[loaf.scala 295:21]
  wire [15:0] _T_1904; // @[loaf.scala 295:34]
  wire  _T_1906; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2201; // @[loaf.scala 298:37]
  wire [21:0] _T_1908; // @[loaf.scala 316:29]
  wire  _T_1910; // @[loaf.scala 292:22]
  wire [15:0] _T_1912; // @[loaf.scala 294:33]
  wire  _T_1914; // @[loaf.scala 295:21]
  wire [15:0] _T_1916; // @[loaf.scala 295:34]
  wire  _T_1918; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2204; // @[loaf.scala 298:37]
  wire [21:0] _T_1920; // @[loaf.scala 316:29]
  wire  _T_1922; // @[loaf.scala 292:22]
  wire [15:0] _T_1924; // @[loaf.scala 294:33]
  wire  _T_1926; // @[loaf.scala 295:21]
  wire [15:0] _T_1928; // @[loaf.scala 295:34]
  wire  _T_1930; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2207; // @[loaf.scala 298:37]
  wire [21:0] _T_1932; // @[loaf.scala 316:29]
  wire  _T_1934; // @[loaf.scala 292:22]
  wire [15:0] _T_1936; // @[loaf.scala 294:33]
  wire  _T_1938; // @[loaf.scala 295:21]
  wire [15:0] _T_1940; // @[loaf.scala 295:34]
  wire  _T_1942; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2210; // @[loaf.scala 298:37]
  wire [21:0] _T_1944; // @[loaf.scala 316:29]
  wire  _T_1946; // @[loaf.scala 292:22]
  wire [15:0] _T_1948; // @[loaf.scala 294:33]
  wire  _T_1950; // @[loaf.scala 295:21]
  wire [15:0] _T_1952; // @[loaf.scala 295:34]
  wire  _T_1954; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2213; // @[loaf.scala 298:37]
  wire [21:0] _T_1956; // @[loaf.scala 316:29]
  wire  _T_1958; // @[loaf.scala 292:22]
  wire [15:0] _T_1960; // @[loaf.scala 294:33]
  wire  _T_1962; // @[loaf.scala 295:21]
  wire [15:0] _T_1964; // @[loaf.scala 295:34]
  wire  _T_1966; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2216; // @[loaf.scala 298:37]
  wire [21:0] _T_1968; // @[loaf.scala 316:29]
  wire  _T_1970; // @[loaf.scala 327:24]
  wire [21:0] _GEN_2217; // @[loaf.scala 327:29]
  wire  _T_1972; // @[loaf.scala 327:24]
  wire [21:0] _GEN_2218; // @[loaf.scala 327:29]
  wire  _T_1974; // @[loaf.scala 327:24]
  wire [21:0] _GEN_2219; // @[loaf.scala 327:29]
  wire  _T_1976; // @[loaf.scala 327:24]
  wire [21:0] _GEN_2220; // @[loaf.scala 327:29]
  wire  _T_1978; // @[loaf.scala 327:24]
  wire  _T_1980; // @[loaf.scala 327:24]
  wire  _T_1982; // @[loaf.scala 327:24]
  wire  _T_1984; // @[loaf.scala 354:43]
  wire  _T_1985; // @[loaf.scala 354:35]
  wire  _T_1987; // @[loaf.scala 292:22]
  wire [15:0] _T_1989; // @[loaf.scala 294:33]
  wire  _T_1991; // @[loaf.scala 295:21]
  wire [15:0] _T_1993; // @[loaf.scala 295:34]
  wire  _T_1995; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2227; // @[loaf.scala 298:37]
  wire [21:0] _T_1997; // @[loaf.scala 316:29]
  wire  _T_1999; // @[loaf.scala 292:22]
  wire [15:0] _T_2001; // @[loaf.scala 294:33]
  wire  _T_2003; // @[loaf.scala 295:21]
  wire [15:0] _T_2005; // @[loaf.scala 295:34]
  wire  _T_2007; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2230; // @[loaf.scala 298:37]
  wire [21:0] _T_2009; // @[loaf.scala 316:29]
  wire  _T_2011; // @[loaf.scala 292:22]
  wire [15:0] _T_2013; // @[loaf.scala 294:33]
  wire  _T_2015; // @[loaf.scala 295:21]
  wire [15:0] _T_2017; // @[loaf.scala 295:34]
  wire  _T_2019; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2233; // @[loaf.scala 298:37]
  wire [21:0] _T_2021; // @[loaf.scala 316:29]
  wire  _T_2023; // @[loaf.scala 292:22]
  wire [15:0] _T_2025; // @[loaf.scala 294:33]
  wire  _T_2027; // @[loaf.scala 295:21]
  wire [15:0] _T_2029; // @[loaf.scala 295:34]
  wire  _T_2031; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2236; // @[loaf.scala 298:37]
  wire [21:0] _T_2033; // @[loaf.scala 316:29]
  wire  _T_2035; // @[loaf.scala 292:22]
  wire [15:0] _T_2037; // @[loaf.scala 294:33]
  wire  _T_2039; // @[loaf.scala 295:21]
  wire [15:0] _T_2041; // @[loaf.scala 295:34]
  wire  _T_2043; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2239; // @[loaf.scala 298:37]
  wire [21:0] _T_2045; // @[loaf.scala 316:29]
  wire  _T_2047; // @[loaf.scala 292:22]
  wire [15:0] _T_2049; // @[loaf.scala 294:33]
  wire  _T_2051; // @[loaf.scala 295:21]
  wire [15:0] _T_2053; // @[loaf.scala 295:34]
  wire  _T_2055; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2242; // @[loaf.scala 298:37]
  wire [21:0] _T_2057; // @[loaf.scala 316:29]
  wire  _T_2059; // @[loaf.scala 292:22]
  wire [15:0] _T_2061; // @[loaf.scala 294:33]
  wire  _T_2063; // @[loaf.scala 295:21]
  wire [15:0] _T_2065; // @[loaf.scala 295:34]
  wire  _T_2067; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2245; // @[loaf.scala 298:37]
  wire [21:0] _T_2069; // @[loaf.scala 316:29]
  wire  _T_2071; // @[loaf.scala 292:22]
  wire [15:0] _T_2073; // @[loaf.scala 294:33]
  wire  _T_2075; // @[loaf.scala 295:21]
  wire [15:0] _T_2077; // @[loaf.scala 295:34]
  wire  _T_2079; // @[loaf.scala 298:29]
  wire [15:0] _GEN_2248; // @[loaf.scala 298:37]
  wire [21:0] _T_2081; // @[loaf.scala 316:29]
  wire  _T_2083; // @[loaf.scala 327:24]
  wire [21:0] _GEN_2249; // @[loaf.scala 327:29]
  wire  _T_2085; // @[loaf.scala 327:24]
  wire [21:0] _GEN_2250; // @[loaf.scala 327:29]
  wire  _T_2087; // @[loaf.scala 327:24]
  wire [21:0] _GEN_2251; // @[loaf.scala 327:29]
  wire  _T_2089; // @[loaf.scala 327:24]
  wire [21:0] _GEN_2252; // @[loaf.scala 327:29]
  wire  _T_2091; // @[loaf.scala 327:24]
  wire  _T_2093; // @[loaf.scala 327:24]
  wire  _T_2095; // @[loaf.scala 327:24]
  wire  _T_2097; // @[loaf.scala 354:43]
  wire  _T_2098; // @[loaf.scala 354:35]
  wire  _T_2102; // @[loaf.scala 363:20]
  wire [1:0] _T_2104; // @[loaf.scala 364:20]
  wire  _T_2105; // @[loaf.scala 367:22]
  wire [1:0] _T_2107; // @[loaf.scala 368:22]
  wire  _T_2108; // @[loaf.scala 375:31]
  wire [8:0] _T_2110; // @[loaf.scala 376:36]
  wire  _T_2112; // @[loaf.scala 388:75]
  wire  _T_2114; // @[loaf.scala 388:75]
  wire  _T_2115; // @[loaf.scala 388:72]
  wire  _T_2116; // @[loaf.scala 388:75]
  wire  _T_2117; // @[loaf.scala 388:72]
  wire  _T_2118; // @[loaf.scala 388:75]
  wire  _T_2119; // @[loaf.scala 388:72]
  wire  _T_2120; // @[loaf.scala 388:75]
  wire  _T_2121; // @[loaf.scala 388:72]
  wire  _T_2122; // @[loaf.scala 388:75]
  wire  _T_2123; // @[loaf.scala 388:72]
  wire  _T_2124; // @[loaf.scala 388:75]
  wire  _T_2125; // @[loaf.scala 388:72]
  wire  _T_2126; // @[loaf.scala 388:75]
  wire  _T_2127; // @[loaf.scala 388:72]
  wire  _T_2128; // @[loaf.scala 388:75]
  wire  _T_2129; // @[loaf.scala 388:72]
  wire  _T_2130; // @[loaf.scala 388:75]
  wire  _T_2131; // @[loaf.scala 388:72]
  wire  _T_2132; // @[loaf.scala 388:75]
  wire  _T_2133; // @[loaf.scala 388:72]
  wire  _T_2134; // @[loaf.scala 388:75]
  wire  _T_2135; // @[loaf.scala 388:72]
  wire  _T_2136; // @[loaf.scala 388:75]
  wire  _T_2137; // @[loaf.scala 388:72]
  wire  _T_2138; // @[loaf.scala 388:75]
  wire  _T_2139; // @[loaf.scala 388:72]
  wire  _GEN_2323; // @[loaf.scala 246:49]
  wire  _GEN_2324; // @[loaf.scala 246:49]
  wire  _GEN_2365; // @[loaf.scala 246:49]
  wire  _GEN_2370; // @[loaf.scala 246:49]
  wire [25:0] _GEN_2573; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2574; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2575; // @[loaf.scala 246:49]
  wire [25:0] _GEN_2578; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2579; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2580; // @[loaf.scala 246:49]
  wire [25:0] _GEN_2583; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2584; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2585; // @[loaf.scala 246:49]
  wire [25:0] _GEN_2588; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2589; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2590; // @[loaf.scala 246:49]
  wire [25:0] _GEN_2593; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2594; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2595; // @[loaf.scala 246:49]
  wire [25:0] _GEN_2598; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2599; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2600; // @[loaf.scala 246:49]
  wire [25:0] _GEN_2603; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2604; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2605; // @[loaf.scala 246:49]
  wire [25:0] _GEN_2608; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2609; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2610; // @[loaf.scala 246:49]
  wire [21:0] _GEN_2611; // @[loaf.scala 246:49]
  wire [21:0] _GEN_2612; // @[loaf.scala 246:49]
  wire [21:0] _GEN_2613; // @[loaf.scala 246:49]
  wire [21:0] _GEN_2614; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2624; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2625; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2629; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2630; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2634; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2635; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2639; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2640; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2644; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2645; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2649; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2650; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2654; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2655; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2659; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2660; // @[loaf.scala 246:49]
  wire [21:0] _GEN_2661; // @[loaf.scala 246:49]
  wire [21:0] _GEN_2662; // @[loaf.scala 246:49]
  wire [21:0] _GEN_2663; // @[loaf.scala 246:49]
  wire [21:0] _GEN_2664; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2674; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2675; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2679; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2680; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2684; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2685; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2689; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2690; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2694; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2695; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2699; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2700; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2704; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2705; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2709; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2710; // @[loaf.scala 246:49]
  wire [21:0] _GEN_2711; // @[loaf.scala 246:49]
  wire [21:0] _GEN_2712; // @[loaf.scala 246:49]
  wire [21:0] _GEN_2713; // @[loaf.scala 246:49]
  wire [21:0] _GEN_2714; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2724; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2725; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2729; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2730; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2734; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2735; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2739; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2740; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2744; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2745; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2749; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2750; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2754; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2755; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2759; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2760; // @[loaf.scala 246:49]
  wire [21:0] _GEN_2761; // @[loaf.scala 246:49]
  wire [21:0] _GEN_2762; // @[loaf.scala 246:49]
  wire [21:0] _GEN_2763; // @[loaf.scala 246:49]
  wire [21:0] _GEN_2764; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2774; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2775; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2779; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2780; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2784; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2785; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2789; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2790; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2794; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2795; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2799; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2800; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2804; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2805; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2809; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2810; // @[loaf.scala 246:49]
  wire [21:0] _GEN_2811; // @[loaf.scala 246:49]
  wire [21:0] _GEN_2812; // @[loaf.scala 246:49]
  wire [21:0] _GEN_2813; // @[loaf.scala 246:49]
  wire [21:0] _GEN_2814; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2824; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2825; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2829; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2830; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2834; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2835; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2839; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2840; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2844; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2845; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2849; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2850; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2854; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2855; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2859; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2860; // @[loaf.scala 246:49]
  wire [21:0] _GEN_2861; // @[loaf.scala 246:49]
  wire [21:0] _GEN_2862; // @[loaf.scala 246:49]
  wire [21:0] _GEN_2863; // @[loaf.scala 246:49]
  wire [21:0] _GEN_2864; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2874; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2875; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2879; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2880; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2884; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2885; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2889; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2890; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2894; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2895; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2899; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2900; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2904; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2905; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2909; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2910; // @[loaf.scala 246:49]
  wire [21:0] _GEN_2911; // @[loaf.scala 246:49]
  wire [21:0] _GEN_2912; // @[loaf.scala 246:49]
  wire [21:0] _GEN_2913; // @[loaf.scala 246:49]
  wire [21:0] _GEN_2914; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2924; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2925; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2929; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2930; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2934; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2935; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2939; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2940; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2944; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2945; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2949; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2950; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2954; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2955; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2959; // @[loaf.scala 246:49]
  wire [15:0] _GEN_2960; // @[loaf.scala 246:49]
  wire [21:0] _GEN_2961; // @[loaf.scala 246:49]
  wire [21:0] _GEN_2962; // @[loaf.scala 246:49]
  wire [21:0] _GEN_2963; // @[loaf.scala 246:49]
  wire [21:0] _GEN_2964; // @[loaf.scala 246:49]
  wire  _GEN_3036; // @[loaf.scala 236:43]
  wire  _GEN_3037; // @[loaf.scala 236:43]
  wire  _GEN_3078; // @[loaf.scala 236:43]
  wire  _GEN_3083; // @[loaf.scala 236:43]
  wire  _GEN_3285; // @[loaf.scala 236:43]
  wire [25:0] _GEN_3286; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3287; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3288; // @[loaf.scala 236:43]
  wire [25:0] _GEN_3291; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3292; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3293; // @[loaf.scala 236:43]
  wire [25:0] _GEN_3296; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3297; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3298; // @[loaf.scala 236:43]
  wire [25:0] _GEN_3301; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3302; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3303; // @[loaf.scala 236:43]
  wire [25:0] _GEN_3306; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3307; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3308; // @[loaf.scala 236:43]
  wire [25:0] _GEN_3311; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3312; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3313; // @[loaf.scala 236:43]
  wire [25:0] _GEN_3316; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3317; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3318; // @[loaf.scala 236:43]
  wire [25:0] _GEN_3321; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3322; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3323; // @[loaf.scala 236:43]
  wire [21:0] _GEN_3324; // @[loaf.scala 236:43]
  wire [21:0] _GEN_3325; // @[loaf.scala 236:43]
  wire [21:0] _GEN_3326; // @[loaf.scala 236:43]
  wire [21:0] _GEN_3327; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3337; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3338; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3342; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3343; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3347; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3348; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3352; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3353; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3357; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3358; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3362; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3363; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3367; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3368; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3372; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3373; // @[loaf.scala 236:43]
  wire [21:0] _GEN_3374; // @[loaf.scala 236:43]
  wire [21:0] _GEN_3375; // @[loaf.scala 236:43]
  wire [21:0] _GEN_3376; // @[loaf.scala 236:43]
  wire [21:0] _GEN_3377; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3387; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3388; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3392; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3393; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3397; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3398; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3402; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3403; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3407; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3408; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3412; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3413; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3417; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3418; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3422; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3423; // @[loaf.scala 236:43]
  wire [21:0] _GEN_3424; // @[loaf.scala 236:43]
  wire [21:0] _GEN_3425; // @[loaf.scala 236:43]
  wire [21:0] _GEN_3426; // @[loaf.scala 236:43]
  wire [21:0] _GEN_3427; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3437; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3438; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3442; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3443; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3447; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3448; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3452; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3453; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3457; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3458; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3462; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3463; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3467; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3468; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3472; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3473; // @[loaf.scala 236:43]
  wire [21:0] _GEN_3474; // @[loaf.scala 236:43]
  wire [21:0] _GEN_3475; // @[loaf.scala 236:43]
  wire [21:0] _GEN_3476; // @[loaf.scala 236:43]
  wire [21:0] _GEN_3477; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3487; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3488; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3492; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3493; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3497; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3498; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3502; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3503; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3507; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3508; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3512; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3513; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3517; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3518; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3522; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3523; // @[loaf.scala 236:43]
  wire [21:0] _GEN_3524; // @[loaf.scala 236:43]
  wire [21:0] _GEN_3525; // @[loaf.scala 236:43]
  wire [21:0] _GEN_3526; // @[loaf.scala 236:43]
  wire [21:0] _GEN_3527; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3537; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3538; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3542; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3543; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3547; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3548; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3552; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3553; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3557; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3558; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3562; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3563; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3567; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3568; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3572; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3573; // @[loaf.scala 236:43]
  wire [21:0] _GEN_3574; // @[loaf.scala 236:43]
  wire [21:0] _GEN_3575; // @[loaf.scala 236:43]
  wire [21:0] _GEN_3576; // @[loaf.scala 236:43]
  wire [21:0] _GEN_3577; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3587; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3588; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3592; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3593; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3597; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3598; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3602; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3603; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3607; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3608; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3612; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3613; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3617; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3618; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3622; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3623; // @[loaf.scala 236:43]
  wire [21:0] _GEN_3624; // @[loaf.scala 236:43]
  wire [21:0] _GEN_3625; // @[loaf.scala 236:43]
  wire [21:0] _GEN_3626; // @[loaf.scala 236:43]
  wire [21:0] _GEN_3627; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3637; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3638; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3642; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3643; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3647; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3648; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3652; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3653; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3657; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3658; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3662; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3663; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3667; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3668; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3672; // @[loaf.scala 236:43]
  wire [15:0] _GEN_3673; // @[loaf.scala 236:43]
  wire [21:0] _GEN_3674; // @[loaf.scala 236:43]
  wire [21:0] _GEN_3675; // @[loaf.scala 236:43]
  wire [21:0] _GEN_3676; // @[loaf.scala 236:43]
  wire [21:0] _GEN_3677; // @[loaf.scala 236:43]
  wire [25:0] _GEN_3998; // @[loaf.scala 234:29]
  wire [25:0] _GEN_4003; // @[loaf.scala 234:29]
  wire [25:0] _GEN_4008; // @[loaf.scala 234:29]
  wire [25:0] _GEN_4013; // @[loaf.scala 234:29]
  wire [25:0] _GEN_4018; // @[loaf.scala 234:29]
  wire [25:0] _GEN_4023; // @[loaf.scala 234:29]
  wire [25:0] _GEN_4028; // @[loaf.scala 234:29]
  wire [25:0] _GEN_4033; // @[loaf.scala 234:29]
  wire [21:0] _GEN_4036; // @[loaf.scala 234:29]
  wire [21:0] _GEN_4037; // @[loaf.scala 234:29]
  wire [21:0] _GEN_4038; // @[loaf.scala 234:29]
  wire [21:0] _GEN_4039; // @[loaf.scala 234:29]
  wire [21:0] _GEN_4086; // @[loaf.scala 234:29]
  wire [21:0] _GEN_4087; // @[loaf.scala 234:29]
  wire [21:0] _GEN_4088; // @[loaf.scala 234:29]
  wire [21:0] _GEN_4089; // @[loaf.scala 234:29]
  wire [21:0] _GEN_4136; // @[loaf.scala 234:29]
  wire [21:0] _GEN_4137; // @[loaf.scala 234:29]
  wire [21:0] _GEN_4138; // @[loaf.scala 234:29]
  wire [21:0] _GEN_4139; // @[loaf.scala 234:29]
  wire [21:0] _GEN_4186; // @[loaf.scala 234:29]
  wire [21:0] _GEN_4187; // @[loaf.scala 234:29]
  wire [21:0] _GEN_4188; // @[loaf.scala 234:29]
  wire [21:0] _GEN_4189; // @[loaf.scala 234:29]
  wire [21:0] _GEN_4236; // @[loaf.scala 234:29]
  wire [21:0] _GEN_4237; // @[loaf.scala 234:29]
  wire [21:0] _GEN_4238; // @[loaf.scala 234:29]
  wire [21:0] _GEN_4239; // @[loaf.scala 234:29]
  wire [21:0] _GEN_4286; // @[loaf.scala 234:29]
  wire [21:0] _GEN_4287; // @[loaf.scala 234:29]
  wire [21:0] _GEN_4288; // @[loaf.scala 234:29]
  wire [21:0] _GEN_4289; // @[loaf.scala 234:29]
  wire [21:0] _GEN_4336; // @[loaf.scala 234:29]
  wire [21:0] _GEN_4337; // @[loaf.scala 234:29]
  wire [21:0] _GEN_4338; // @[loaf.scala 234:29]
  wire [21:0] _GEN_4339; // @[loaf.scala 234:29]
  wire [21:0] _GEN_4386; // @[loaf.scala 234:29]
  wire [21:0] _GEN_4387; // @[loaf.scala 234:29]
  wire [21:0] _GEN_4388; // @[loaf.scala 234:29]
  wire [21:0] _GEN_4389; // @[loaf.scala 234:29]
  wire [15:0] _GEN_4987; // @[loaf.scala 337:25]
  wire [15:0] _GEN_4988; // @[loaf.scala 337:25]
  wire [15:0] _GEN_4989; // @[loaf.scala 337:25]
  wire [15:0] _GEN_4990; // @[loaf.scala 337:25]
  wire [15:0] _GEN_4991; // @[loaf.scala 337:25]
  wire [15:0] _GEN_4992; // @[loaf.scala 337:25]
  wire [15:0] _GEN_4993; // @[loaf.scala 337:25]
  wire [15:0] _GEN_4994; // @[loaf.scala 337:25]
  wire [15:0] _GEN_4995; // @[loaf.scala 337:25]
  wire [15:0] _GEN_4996; // @[loaf.scala 337:25]
  wire [15:0] _GEN_4997; // @[loaf.scala 337:25]
  wire [15:0] _GEN_4998; // @[loaf.scala 337:25]
  wire [15:0] _GEN_4999; // @[loaf.scala 337:25]
  wire [15:0] _GEN_5000; // @[loaf.scala 337:25]
  wire [15:0] _GEN_5001; // @[loaf.scala 337:25]
  wire [15:0] _GEN_5002; // @[loaf.scala 337:25]
  wire [15:0] _GEN_5003; // @[loaf.scala 337:25]
  wire [15:0] _GEN_5004; // @[loaf.scala 337:25]
  wire [15:0] _GEN_5005; // @[loaf.scala 337:25]
  wire [15:0] _GEN_5006; // @[loaf.scala 337:25]
  wire [15:0] _GEN_5007; // @[loaf.scala 337:25]
  wire [15:0] _GEN_5008; // @[loaf.scala 337:25]
  wire [15:0] _GEN_5009; // @[loaf.scala 337:25]
  wire [15:0] _GEN_5010; // @[loaf.scala 337:25]
  wire [15:0] _GEN_5011; // @[loaf.scala 337:25]
  wire [15:0] _GEN_5012; // @[loaf.scala 337:25]
  wire [15:0] _GEN_5013; // @[loaf.scala 337:25]
  wire [15:0] _GEN_5014; // @[loaf.scala 337:25]
  wire [15:0] _GEN_5015; // @[loaf.scala 337:25]
  wire [15:0] _GEN_5016; // @[loaf.scala 337:25]
  wire [15:0] _GEN_5017; // @[loaf.scala 337:25]
  wire [15:0] _GEN_5018; // @[loaf.scala 337:25]
  MAC macs_0_0 ( // @[loaf.scala 120:72]
    .clock(macs_0_0_clock),
    .io_en(macs_0_0_io_en),
    .io_a(macs_0_0_io_a),
    .io_b(macs_0_0_io_b),
    .io_o(macs_0_0_io_o),
    .io_r(macs_0_0_io_r)
  );
  MAC macs_0_1 ( // @[loaf.scala 120:72]
    .clock(macs_0_1_clock),
    .io_en(macs_0_1_io_en),
    .io_a(macs_0_1_io_a),
    .io_b(macs_0_1_io_b),
    .io_o(macs_0_1_io_o),
    .io_r(macs_0_1_io_r)
  );
  MAC macs_0_2 ( // @[loaf.scala 120:72]
    .clock(macs_0_2_clock),
    .io_en(macs_0_2_io_en),
    .io_a(macs_0_2_io_a),
    .io_b(macs_0_2_io_b),
    .io_o(macs_0_2_io_o),
    .io_r(macs_0_2_io_r)
  );
  MAC macs_0_3 ( // @[loaf.scala 120:72]
    .clock(macs_0_3_clock),
    .io_en(macs_0_3_io_en),
    .io_a(macs_0_3_io_a),
    .io_b(macs_0_3_io_b),
    .io_o(macs_0_3_io_o),
    .io_r(macs_0_3_io_r)
  );
  MAC macs_0_4 ( // @[loaf.scala 120:72]
    .clock(macs_0_4_clock),
    .io_en(macs_0_4_io_en),
    .io_a(macs_0_4_io_a),
    .io_b(macs_0_4_io_b),
    .io_o(macs_0_4_io_o),
    .io_r(macs_0_4_io_r)
  );
  MAC macs_0_5 ( // @[loaf.scala 120:72]
    .clock(macs_0_5_clock),
    .io_en(macs_0_5_io_en),
    .io_a(macs_0_5_io_a),
    .io_b(macs_0_5_io_b),
    .io_o(macs_0_5_io_o),
    .io_r(macs_0_5_io_r)
  );
  MAC macs_0_6 ( // @[loaf.scala 120:72]
    .clock(macs_0_6_clock),
    .io_en(macs_0_6_io_en),
    .io_a(macs_0_6_io_a),
    .io_b(macs_0_6_io_b),
    .io_o(macs_0_6_io_o),
    .io_r(macs_0_6_io_r)
  );
  MAC macs_0_7 ( // @[loaf.scala 120:72]
    .clock(macs_0_7_clock),
    .io_en(macs_0_7_io_en),
    .io_a(macs_0_7_io_a),
    .io_b(macs_0_7_io_b),
    .io_o(macs_0_7_io_o),
    .io_r(macs_0_7_io_r)
  );
  MAC macs_1_0 ( // @[loaf.scala 120:72]
    .clock(macs_1_0_clock),
    .io_en(macs_1_0_io_en),
    .io_a(macs_1_0_io_a),
    .io_b(macs_1_0_io_b),
    .io_o(macs_1_0_io_o),
    .io_r(macs_1_0_io_r)
  );
  MAC macs_1_1 ( // @[loaf.scala 120:72]
    .clock(macs_1_1_clock),
    .io_en(macs_1_1_io_en),
    .io_a(macs_1_1_io_a),
    .io_b(macs_1_1_io_b),
    .io_o(macs_1_1_io_o),
    .io_r(macs_1_1_io_r)
  );
  MAC macs_1_2 ( // @[loaf.scala 120:72]
    .clock(macs_1_2_clock),
    .io_en(macs_1_2_io_en),
    .io_a(macs_1_2_io_a),
    .io_b(macs_1_2_io_b),
    .io_o(macs_1_2_io_o),
    .io_r(macs_1_2_io_r)
  );
  MAC macs_1_3 ( // @[loaf.scala 120:72]
    .clock(macs_1_3_clock),
    .io_en(macs_1_3_io_en),
    .io_a(macs_1_3_io_a),
    .io_b(macs_1_3_io_b),
    .io_o(macs_1_3_io_o),
    .io_r(macs_1_3_io_r)
  );
  MAC macs_1_4 ( // @[loaf.scala 120:72]
    .clock(macs_1_4_clock),
    .io_en(macs_1_4_io_en),
    .io_a(macs_1_4_io_a),
    .io_b(macs_1_4_io_b),
    .io_o(macs_1_4_io_o),
    .io_r(macs_1_4_io_r)
  );
  MAC macs_1_5 ( // @[loaf.scala 120:72]
    .clock(macs_1_5_clock),
    .io_en(macs_1_5_io_en),
    .io_a(macs_1_5_io_a),
    .io_b(macs_1_5_io_b),
    .io_o(macs_1_5_io_o),
    .io_r(macs_1_5_io_r)
  );
  MAC macs_1_6 ( // @[loaf.scala 120:72]
    .clock(macs_1_6_clock),
    .io_en(macs_1_6_io_en),
    .io_a(macs_1_6_io_a),
    .io_b(macs_1_6_io_b),
    .io_o(macs_1_6_io_o),
    .io_r(macs_1_6_io_r)
  );
  MAC macs_1_7 ( // @[loaf.scala 120:72]
    .clock(macs_1_7_clock),
    .io_en(macs_1_7_io_en),
    .io_a(macs_1_7_io_a),
    .io_b(macs_1_7_io_b),
    .io_o(macs_1_7_io_o),
    .io_r(macs_1_7_io_r)
  );
  MAC macs_2_0 ( // @[loaf.scala 120:72]
    .clock(macs_2_0_clock),
    .io_en(macs_2_0_io_en),
    .io_a(macs_2_0_io_a),
    .io_b(macs_2_0_io_b),
    .io_o(macs_2_0_io_o),
    .io_r(macs_2_0_io_r)
  );
  MAC macs_2_1 ( // @[loaf.scala 120:72]
    .clock(macs_2_1_clock),
    .io_en(macs_2_1_io_en),
    .io_a(macs_2_1_io_a),
    .io_b(macs_2_1_io_b),
    .io_o(macs_2_1_io_o),
    .io_r(macs_2_1_io_r)
  );
  MAC macs_2_2 ( // @[loaf.scala 120:72]
    .clock(macs_2_2_clock),
    .io_en(macs_2_2_io_en),
    .io_a(macs_2_2_io_a),
    .io_b(macs_2_2_io_b),
    .io_o(macs_2_2_io_o),
    .io_r(macs_2_2_io_r)
  );
  MAC macs_2_3 ( // @[loaf.scala 120:72]
    .clock(macs_2_3_clock),
    .io_en(macs_2_3_io_en),
    .io_a(macs_2_3_io_a),
    .io_b(macs_2_3_io_b),
    .io_o(macs_2_3_io_o),
    .io_r(macs_2_3_io_r)
  );
  MAC macs_2_4 ( // @[loaf.scala 120:72]
    .clock(macs_2_4_clock),
    .io_en(macs_2_4_io_en),
    .io_a(macs_2_4_io_a),
    .io_b(macs_2_4_io_b),
    .io_o(macs_2_4_io_o),
    .io_r(macs_2_4_io_r)
  );
  MAC macs_2_5 ( // @[loaf.scala 120:72]
    .clock(macs_2_5_clock),
    .io_en(macs_2_5_io_en),
    .io_a(macs_2_5_io_a),
    .io_b(macs_2_5_io_b),
    .io_o(macs_2_5_io_o),
    .io_r(macs_2_5_io_r)
  );
  MAC macs_2_6 ( // @[loaf.scala 120:72]
    .clock(macs_2_6_clock),
    .io_en(macs_2_6_io_en),
    .io_a(macs_2_6_io_a),
    .io_b(macs_2_6_io_b),
    .io_o(macs_2_6_io_o),
    .io_r(macs_2_6_io_r)
  );
  MAC macs_2_7 ( // @[loaf.scala 120:72]
    .clock(macs_2_7_clock),
    .io_en(macs_2_7_io_en),
    .io_a(macs_2_7_io_a),
    .io_b(macs_2_7_io_b),
    .io_o(macs_2_7_io_o),
    .io_r(macs_2_7_io_r)
  );
  MAC macs_3_0 ( // @[loaf.scala 120:72]
    .clock(macs_3_0_clock),
    .io_en(macs_3_0_io_en),
    .io_a(macs_3_0_io_a),
    .io_b(macs_3_0_io_b),
    .io_o(macs_3_0_io_o),
    .io_r(macs_3_0_io_r)
  );
  MAC macs_3_1 ( // @[loaf.scala 120:72]
    .clock(macs_3_1_clock),
    .io_en(macs_3_1_io_en),
    .io_a(macs_3_1_io_a),
    .io_b(macs_3_1_io_b),
    .io_o(macs_3_1_io_o),
    .io_r(macs_3_1_io_r)
  );
  MAC macs_3_2 ( // @[loaf.scala 120:72]
    .clock(macs_3_2_clock),
    .io_en(macs_3_2_io_en),
    .io_a(macs_3_2_io_a),
    .io_b(macs_3_2_io_b),
    .io_o(macs_3_2_io_o),
    .io_r(macs_3_2_io_r)
  );
  MAC macs_3_3 ( // @[loaf.scala 120:72]
    .clock(macs_3_3_clock),
    .io_en(macs_3_3_io_en),
    .io_a(macs_3_3_io_a),
    .io_b(macs_3_3_io_b),
    .io_o(macs_3_3_io_o),
    .io_r(macs_3_3_io_r)
  );
  MAC macs_3_4 ( // @[loaf.scala 120:72]
    .clock(macs_3_4_clock),
    .io_en(macs_3_4_io_en),
    .io_a(macs_3_4_io_a),
    .io_b(macs_3_4_io_b),
    .io_o(macs_3_4_io_o),
    .io_r(macs_3_4_io_r)
  );
  MAC macs_3_5 ( // @[loaf.scala 120:72]
    .clock(macs_3_5_clock),
    .io_en(macs_3_5_io_en),
    .io_a(macs_3_5_io_a),
    .io_b(macs_3_5_io_b),
    .io_o(macs_3_5_io_o),
    .io_r(macs_3_5_io_r)
  );
  MAC macs_3_6 ( // @[loaf.scala 120:72]
    .clock(macs_3_6_clock),
    .io_en(macs_3_6_io_en),
    .io_a(macs_3_6_io_a),
    .io_b(macs_3_6_io_b),
    .io_o(macs_3_6_io_o),
    .io_r(macs_3_6_io_r)
  );
  MAC macs_3_7 ( // @[loaf.scala 120:72]
    .clock(macs_3_7_clock),
    .io_en(macs_3_7_io_en),
    .io_a(macs_3_7_io_a),
    .io_b(macs_3_7_io_b),
    .io_o(macs_3_7_io_o),
    .io_r(macs_3_7_io_r)
  );
  MAC macs_4_0 ( // @[loaf.scala 120:72]
    .clock(macs_4_0_clock),
    .io_en(macs_4_0_io_en),
    .io_a(macs_4_0_io_a),
    .io_b(macs_4_0_io_b),
    .io_o(macs_4_0_io_o),
    .io_r(macs_4_0_io_r)
  );
  MAC macs_4_1 ( // @[loaf.scala 120:72]
    .clock(macs_4_1_clock),
    .io_en(macs_4_1_io_en),
    .io_a(macs_4_1_io_a),
    .io_b(macs_4_1_io_b),
    .io_o(macs_4_1_io_o),
    .io_r(macs_4_1_io_r)
  );
  MAC macs_4_2 ( // @[loaf.scala 120:72]
    .clock(macs_4_2_clock),
    .io_en(macs_4_2_io_en),
    .io_a(macs_4_2_io_a),
    .io_b(macs_4_2_io_b),
    .io_o(macs_4_2_io_o),
    .io_r(macs_4_2_io_r)
  );
  MAC macs_4_3 ( // @[loaf.scala 120:72]
    .clock(macs_4_3_clock),
    .io_en(macs_4_3_io_en),
    .io_a(macs_4_3_io_a),
    .io_b(macs_4_3_io_b),
    .io_o(macs_4_3_io_o),
    .io_r(macs_4_3_io_r)
  );
  MAC macs_4_4 ( // @[loaf.scala 120:72]
    .clock(macs_4_4_clock),
    .io_en(macs_4_4_io_en),
    .io_a(macs_4_4_io_a),
    .io_b(macs_4_4_io_b),
    .io_o(macs_4_4_io_o),
    .io_r(macs_4_4_io_r)
  );
  MAC macs_4_5 ( // @[loaf.scala 120:72]
    .clock(macs_4_5_clock),
    .io_en(macs_4_5_io_en),
    .io_a(macs_4_5_io_a),
    .io_b(macs_4_5_io_b),
    .io_o(macs_4_5_io_o),
    .io_r(macs_4_5_io_r)
  );
  MAC macs_4_6 ( // @[loaf.scala 120:72]
    .clock(macs_4_6_clock),
    .io_en(macs_4_6_io_en),
    .io_a(macs_4_6_io_a),
    .io_b(macs_4_6_io_b),
    .io_o(macs_4_6_io_o),
    .io_r(macs_4_6_io_r)
  );
  MAC macs_4_7 ( // @[loaf.scala 120:72]
    .clock(macs_4_7_clock),
    .io_en(macs_4_7_io_en),
    .io_a(macs_4_7_io_a),
    .io_b(macs_4_7_io_b),
    .io_o(macs_4_7_io_o),
    .io_r(macs_4_7_io_r)
  );
  MAC macs_5_0 ( // @[loaf.scala 120:72]
    .clock(macs_5_0_clock),
    .io_en(macs_5_0_io_en),
    .io_a(macs_5_0_io_a),
    .io_b(macs_5_0_io_b),
    .io_o(macs_5_0_io_o),
    .io_r(macs_5_0_io_r)
  );
  MAC macs_5_1 ( // @[loaf.scala 120:72]
    .clock(macs_5_1_clock),
    .io_en(macs_5_1_io_en),
    .io_a(macs_5_1_io_a),
    .io_b(macs_5_1_io_b),
    .io_o(macs_5_1_io_o),
    .io_r(macs_5_1_io_r)
  );
  MAC macs_5_2 ( // @[loaf.scala 120:72]
    .clock(macs_5_2_clock),
    .io_en(macs_5_2_io_en),
    .io_a(macs_5_2_io_a),
    .io_b(macs_5_2_io_b),
    .io_o(macs_5_2_io_o),
    .io_r(macs_5_2_io_r)
  );
  MAC macs_5_3 ( // @[loaf.scala 120:72]
    .clock(macs_5_3_clock),
    .io_en(macs_5_3_io_en),
    .io_a(macs_5_3_io_a),
    .io_b(macs_5_3_io_b),
    .io_o(macs_5_3_io_o),
    .io_r(macs_5_3_io_r)
  );
  MAC macs_5_4 ( // @[loaf.scala 120:72]
    .clock(macs_5_4_clock),
    .io_en(macs_5_4_io_en),
    .io_a(macs_5_4_io_a),
    .io_b(macs_5_4_io_b),
    .io_o(macs_5_4_io_o),
    .io_r(macs_5_4_io_r)
  );
  MAC macs_5_5 ( // @[loaf.scala 120:72]
    .clock(macs_5_5_clock),
    .io_en(macs_5_5_io_en),
    .io_a(macs_5_5_io_a),
    .io_b(macs_5_5_io_b),
    .io_o(macs_5_5_io_o),
    .io_r(macs_5_5_io_r)
  );
  MAC macs_5_6 ( // @[loaf.scala 120:72]
    .clock(macs_5_6_clock),
    .io_en(macs_5_6_io_en),
    .io_a(macs_5_6_io_a),
    .io_b(macs_5_6_io_b),
    .io_o(macs_5_6_io_o),
    .io_r(macs_5_6_io_r)
  );
  MAC macs_5_7 ( // @[loaf.scala 120:72]
    .clock(macs_5_7_clock),
    .io_en(macs_5_7_io_en),
    .io_a(macs_5_7_io_a),
    .io_b(macs_5_7_io_b),
    .io_o(macs_5_7_io_o),
    .io_r(macs_5_7_io_r)
  );
  MAC macs_6_0 ( // @[loaf.scala 120:72]
    .clock(macs_6_0_clock),
    .io_en(macs_6_0_io_en),
    .io_a(macs_6_0_io_a),
    .io_b(macs_6_0_io_b),
    .io_o(macs_6_0_io_o),
    .io_r(macs_6_0_io_r)
  );
  MAC macs_6_1 ( // @[loaf.scala 120:72]
    .clock(macs_6_1_clock),
    .io_en(macs_6_1_io_en),
    .io_a(macs_6_1_io_a),
    .io_b(macs_6_1_io_b),
    .io_o(macs_6_1_io_o),
    .io_r(macs_6_1_io_r)
  );
  MAC macs_6_2 ( // @[loaf.scala 120:72]
    .clock(macs_6_2_clock),
    .io_en(macs_6_2_io_en),
    .io_a(macs_6_2_io_a),
    .io_b(macs_6_2_io_b),
    .io_o(macs_6_2_io_o),
    .io_r(macs_6_2_io_r)
  );
  MAC macs_6_3 ( // @[loaf.scala 120:72]
    .clock(macs_6_3_clock),
    .io_en(macs_6_3_io_en),
    .io_a(macs_6_3_io_a),
    .io_b(macs_6_3_io_b),
    .io_o(macs_6_3_io_o),
    .io_r(macs_6_3_io_r)
  );
  MAC macs_6_4 ( // @[loaf.scala 120:72]
    .clock(macs_6_4_clock),
    .io_en(macs_6_4_io_en),
    .io_a(macs_6_4_io_a),
    .io_b(macs_6_4_io_b),
    .io_o(macs_6_4_io_o),
    .io_r(macs_6_4_io_r)
  );
  MAC macs_6_5 ( // @[loaf.scala 120:72]
    .clock(macs_6_5_clock),
    .io_en(macs_6_5_io_en),
    .io_a(macs_6_5_io_a),
    .io_b(macs_6_5_io_b),
    .io_o(macs_6_5_io_o),
    .io_r(macs_6_5_io_r)
  );
  MAC macs_6_6 ( // @[loaf.scala 120:72]
    .clock(macs_6_6_clock),
    .io_en(macs_6_6_io_en),
    .io_a(macs_6_6_io_a),
    .io_b(macs_6_6_io_b),
    .io_o(macs_6_6_io_o),
    .io_r(macs_6_6_io_r)
  );
  MAC macs_6_7 ( // @[loaf.scala 120:72]
    .clock(macs_6_7_clock),
    .io_en(macs_6_7_io_en),
    .io_a(macs_6_7_io_a),
    .io_b(macs_6_7_io_b),
    .io_o(macs_6_7_io_o),
    .io_r(macs_6_7_io_r)
  );
  MAC macs_7_0 ( // @[loaf.scala 120:72]
    .clock(macs_7_0_clock),
    .io_en(macs_7_0_io_en),
    .io_a(macs_7_0_io_a),
    .io_b(macs_7_0_io_b),
    .io_o(macs_7_0_io_o),
    .io_r(macs_7_0_io_r)
  );
  MAC macs_7_1 ( // @[loaf.scala 120:72]
    .clock(macs_7_1_clock),
    .io_en(macs_7_1_io_en),
    .io_a(macs_7_1_io_a),
    .io_b(macs_7_1_io_b),
    .io_o(macs_7_1_io_o),
    .io_r(macs_7_1_io_r)
  );
  MAC macs_7_2 ( // @[loaf.scala 120:72]
    .clock(macs_7_2_clock),
    .io_en(macs_7_2_io_en),
    .io_a(macs_7_2_io_a),
    .io_b(macs_7_2_io_b),
    .io_o(macs_7_2_io_o),
    .io_r(macs_7_2_io_r)
  );
  MAC macs_7_3 ( // @[loaf.scala 120:72]
    .clock(macs_7_3_clock),
    .io_en(macs_7_3_io_en),
    .io_a(macs_7_3_io_a),
    .io_b(macs_7_3_io_b),
    .io_o(macs_7_3_io_o),
    .io_r(macs_7_3_io_r)
  );
  MAC macs_7_4 ( // @[loaf.scala 120:72]
    .clock(macs_7_4_clock),
    .io_en(macs_7_4_io_en),
    .io_a(macs_7_4_io_a),
    .io_b(macs_7_4_io_b),
    .io_o(macs_7_4_io_o),
    .io_r(macs_7_4_io_r)
  );
  MAC macs_7_5 ( // @[loaf.scala 120:72]
    .clock(macs_7_5_clock),
    .io_en(macs_7_5_io_en),
    .io_a(macs_7_5_io_a),
    .io_b(macs_7_5_io_b),
    .io_o(macs_7_5_io_o),
    .io_r(macs_7_5_io_r)
  );
  MAC macs_7_6 ( // @[loaf.scala 120:72]
    .clock(macs_7_6_clock),
    .io_en(macs_7_6_io_en),
    .io_a(macs_7_6_io_a),
    .io_b(macs_7_6_io_b),
    .io_o(macs_7_6_io_o),
    .io_r(macs_7_6_io_r)
  );
  MAC macs_7_7 ( // @[loaf.scala 120:72]
    .clock(macs_7_7_clock),
    .io_en(macs_7_7_io_en),
    .io_a(macs_7_7_io_a),
    .io_b(macs_7_7_io_b),
    .io_o(macs_7_7_io_o),
    .io_r(macs_7_7_io_r)
  );
  assign AE_0_0__T_497_addr = _T_494 + _GEN_4796;
  assign AE_0_0__T_497_data = AE_0_0[AE_0_0__T_497_addr]; // @[loaf.scala 147:67]
  assign AE_0_0__T_9_data = {slcBuf_e,slcBuf_a};
  assign AE_0_0__T_9_addr = prev_idx;
  assign AE_0_0__T_9_mask = 1'h1;
  assign AE_0_0__T_9_en = _T_2 ? _GEN_989 : 1'h0;
  assign AE_0_1__T_585_addr = _T_494 + _GEN_4796;
  assign AE_0_1__T_585_data = AE_0_1[AE_0_1__T_585_addr]; // @[loaf.scala 147:67]
  assign AE_0_1__T_15_data = {slcBuf_e,slcBuf_a};
  assign AE_0_1__T_15_addr = prev_idx;
  assign AE_0_1__T_15_mask = 1'h1;
  assign AE_0_1__T_15_en = _T_2 ? _GEN_994 : 1'h0;
  assign AE_0_2__T_673_addr = _T_494 + _GEN_4796;
  assign AE_0_2__T_673_data = AE_0_2[AE_0_2__T_673_addr]; // @[loaf.scala 147:67]
  assign AE_0_2__T_21_data = {slcBuf_e,slcBuf_a};
  assign AE_0_2__T_21_addr = prev_idx;
  assign AE_0_2__T_21_mask = 1'h1;
  assign AE_0_2__T_21_en = _T_2 ? _GEN_999 : 1'h0;
  assign AE_0_3__T_761_addr = _T_494 + _GEN_4796;
  assign AE_0_3__T_761_data = AE_0_3[AE_0_3__T_761_addr]; // @[loaf.scala 147:67]
  assign AE_0_3__T_27_data = {slcBuf_e,slcBuf_a};
  assign AE_0_3__T_27_addr = prev_idx;
  assign AE_0_3__T_27_mask = 1'h1;
  assign AE_0_3__T_27_en = _T_2 ? _GEN_1004 : 1'h0;
  assign AE_0_4__T_849_addr = _T_494 + _GEN_4796;
  assign AE_0_4__T_849_data = AE_0_4[AE_0_4__T_849_addr]; // @[loaf.scala 147:67]
  assign AE_0_4__T_33_data = {slcBuf_e,slcBuf_a};
  assign AE_0_4__T_33_addr = prev_idx;
  assign AE_0_4__T_33_mask = 1'h1;
  assign AE_0_4__T_33_en = _T_2 ? _GEN_1009 : 1'h0;
  assign AE_0_5__T_937_addr = _T_494 + _GEN_4796;
  assign AE_0_5__T_937_data = AE_0_5[AE_0_5__T_937_addr]; // @[loaf.scala 147:67]
  assign AE_0_5__T_39_data = {slcBuf_e,slcBuf_a};
  assign AE_0_5__T_39_addr = prev_idx;
  assign AE_0_5__T_39_mask = 1'h1;
  assign AE_0_5__T_39_en = _T_2 ? _GEN_1014 : 1'h0;
  assign AE_0_6__T_1025_addr = _T_494 + _GEN_4796;
  assign AE_0_6__T_1025_data = AE_0_6[AE_0_6__T_1025_addr]; // @[loaf.scala 147:67]
  assign AE_0_6__T_45_data = {slcBuf_e,slcBuf_a};
  assign AE_0_6__T_45_addr = prev_idx;
  assign AE_0_6__T_45_mask = 1'h1;
  assign AE_0_6__T_45_en = _T_2 ? _GEN_1019 : 1'h0;
  assign AE_0_7__T_1113_addr = _T_494 + _GEN_4796;
  assign AE_0_7__T_1113_data = AE_0_7[AE_0_7__T_1113_addr]; // @[loaf.scala 147:67]
  assign AE_0_7__T_51_data = {slcBuf_e,slcBuf_a};
  assign AE_0_7__T_51_addr = prev_idx;
  assign AE_0_7__T_51_mask = 1'h1;
  assign AE_0_7__T_51_en = _T_2 ? _GEN_1024 : 1'h0;
  assign AE_1_0__T_508_addr = _T_494 + _GEN_4796;
  assign AE_1_0__T_508_data = AE_1_0[AE_1_0__T_508_addr]; // @[loaf.scala 147:67]
  assign AE_1_0__T_57_data = {slcBuf_e,slcBuf_a};
  assign AE_1_0__T_57_addr = prev_idx;
  assign AE_1_0__T_57_mask = 1'h1;
  assign AE_1_0__T_57_en = _T_2 ? _GEN_1029 : 1'h0;
  assign AE_1_1__T_596_addr = _T_494 + _GEN_4796;
  assign AE_1_1__T_596_data = AE_1_1[AE_1_1__T_596_addr]; // @[loaf.scala 147:67]
  assign AE_1_1__T_63_data = {slcBuf_e,slcBuf_a};
  assign AE_1_1__T_63_addr = prev_idx;
  assign AE_1_1__T_63_mask = 1'h1;
  assign AE_1_1__T_63_en = _T_2 ? _GEN_1034 : 1'h0;
  assign AE_1_2__T_684_addr = _T_494 + _GEN_4796;
  assign AE_1_2__T_684_data = AE_1_2[AE_1_2__T_684_addr]; // @[loaf.scala 147:67]
  assign AE_1_2__T_69_data = {slcBuf_e,slcBuf_a};
  assign AE_1_2__T_69_addr = prev_idx;
  assign AE_1_2__T_69_mask = 1'h1;
  assign AE_1_2__T_69_en = _T_2 ? _GEN_1039 : 1'h0;
  assign AE_1_3__T_772_addr = _T_494 + _GEN_4796;
  assign AE_1_3__T_772_data = AE_1_3[AE_1_3__T_772_addr]; // @[loaf.scala 147:67]
  assign AE_1_3__T_75_data = {slcBuf_e,slcBuf_a};
  assign AE_1_3__T_75_addr = prev_idx;
  assign AE_1_3__T_75_mask = 1'h1;
  assign AE_1_3__T_75_en = _T_2 ? _GEN_1044 : 1'h0;
  assign AE_1_4__T_860_addr = _T_494 + _GEN_4796;
  assign AE_1_4__T_860_data = AE_1_4[AE_1_4__T_860_addr]; // @[loaf.scala 147:67]
  assign AE_1_4__T_81_data = {slcBuf_e,slcBuf_a};
  assign AE_1_4__T_81_addr = prev_idx;
  assign AE_1_4__T_81_mask = 1'h1;
  assign AE_1_4__T_81_en = _T_2 ? _GEN_1049 : 1'h0;
  assign AE_1_5__T_948_addr = _T_494 + _GEN_4796;
  assign AE_1_5__T_948_data = AE_1_5[AE_1_5__T_948_addr]; // @[loaf.scala 147:67]
  assign AE_1_5__T_87_data = {slcBuf_e,slcBuf_a};
  assign AE_1_5__T_87_addr = prev_idx;
  assign AE_1_5__T_87_mask = 1'h1;
  assign AE_1_5__T_87_en = _T_2 ? _GEN_1054 : 1'h0;
  assign AE_1_6__T_1036_addr = _T_494 + _GEN_4796;
  assign AE_1_6__T_1036_data = AE_1_6[AE_1_6__T_1036_addr]; // @[loaf.scala 147:67]
  assign AE_1_6__T_93_data = {slcBuf_e,slcBuf_a};
  assign AE_1_6__T_93_addr = prev_idx;
  assign AE_1_6__T_93_mask = 1'h1;
  assign AE_1_6__T_93_en = _T_2 ? _GEN_1059 : 1'h0;
  assign AE_1_7__T_1124_addr = _T_494 + _GEN_4796;
  assign AE_1_7__T_1124_data = AE_1_7[AE_1_7__T_1124_addr]; // @[loaf.scala 147:67]
  assign AE_1_7__T_99_data = {slcBuf_e,slcBuf_a};
  assign AE_1_7__T_99_addr = prev_idx;
  assign AE_1_7__T_99_mask = 1'h1;
  assign AE_1_7__T_99_en = _T_2 ? _GEN_1064 : 1'h0;
  assign AE_2_0__T_519_addr = _T_494 + _GEN_4796;
  assign AE_2_0__T_519_data = AE_2_0[AE_2_0__T_519_addr]; // @[loaf.scala 147:67]
  assign AE_2_0__T_105_data = {slcBuf_e,slcBuf_a};
  assign AE_2_0__T_105_addr = prev_idx;
  assign AE_2_0__T_105_mask = 1'h1;
  assign AE_2_0__T_105_en = _T_2 ? _GEN_1069 : 1'h0;
  assign AE_2_1__T_607_addr = _T_494 + _GEN_4796;
  assign AE_2_1__T_607_data = AE_2_1[AE_2_1__T_607_addr]; // @[loaf.scala 147:67]
  assign AE_2_1__T_111_data = {slcBuf_e,slcBuf_a};
  assign AE_2_1__T_111_addr = prev_idx;
  assign AE_2_1__T_111_mask = 1'h1;
  assign AE_2_1__T_111_en = _T_2 ? _GEN_1074 : 1'h0;
  assign AE_2_2__T_695_addr = _T_494 + _GEN_4796;
  assign AE_2_2__T_695_data = AE_2_2[AE_2_2__T_695_addr]; // @[loaf.scala 147:67]
  assign AE_2_2__T_117_data = {slcBuf_e,slcBuf_a};
  assign AE_2_2__T_117_addr = prev_idx;
  assign AE_2_2__T_117_mask = 1'h1;
  assign AE_2_2__T_117_en = _T_2 ? _GEN_1079 : 1'h0;
  assign AE_2_3__T_783_addr = _T_494 + _GEN_4796;
  assign AE_2_3__T_783_data = AE_2_3[AE_2_3__T_783_addr]; // @[loaf.scala 147:67]
  assign AE_2_3__T_123_data = {slcBuf_e,slcBuf_a};
  assign AE_2_3__T_123_addr = prev_idx;
  assign AE_2_3__T_123_mask = 1'h1;
  assign AE_2_3__T_123_en = _T_2 ? _GEN_1084 : 1'h0;
  assign AE_2_4__T_871_addr = _T_494 + _GEN_4796;
  assign AE_2_4__T_871_data = AE_2_4[AE_2_4__T_871_addr]; // @[loaf.scala 147:67]
  assign AE_2_4__T_129_data = {slcBuf_e,slcBuf_a};
  assign AE_2_4__T_129_addr = prev_idx;
  assign AE_2_4__T_129_mask = 1'h1;
  assign AE_2_4__T_129_en = _T_2 ? _GEN_1089 : 1'h0;
  assign AE_2_5__T_959_addr = _T_494 + _GEN_4796;
  assign AE_2_5__T_959_data = AE_2_5[AE_2_5__T_959_addr]; // @[loaf.scala 147:67]
  assign AE_2_5__T_135_data = {slcBuf_e,slcBuf_a};
  assign AE_2_5__T_135_addr = prev_idx;
  assign AE_2_5__T_135_mask = 1'h1;
  assign AE_2_5__T_135_en = _T_2 ? _GEN_1094 : 1'h0;
  assign AE_2_6__T_1047_addr = _T_494 + _GEN_4796;
  assign AE_2_6__T_1047_data = AE_2_6[AE_2_6__T_1047_addr]; // @[loaf.scala 147:67]
  assign AE_2_6__T_141_data = {slcBuf_e,slcBuf_a};
  assign AE_2_6__T_141_addr = prev_idx;
  assign AE_2_6__T_141_mask = 1'h1;
  assign AE_2_6__T_141_en = _T_2 ? _GEN_1099 : 1'h0;
  assign AE_2_7__T_1135_addr = _T_494 + _GEN_4796;
  assign AE_2_7__T_1135_data = AE_2_7[AE_2_7__T_1135_addr]; // @[loaf.scala 147:67]
  assign AE_2_7__T_147_data = {slcBuf_e,slcBuf_a};
  assign AE_2_7__T_147_addr = prev_idx;
  assign AE_2_7__T_147_mask = 1'h1;
  assign AE_2_7__T_147_en = _T_2 ? _GEN_1104 : 1'h0;
  assign AE_3_0__T_530_addr = _T_494 + _GEN_4796;
  assign AE_3_0__T_530_data = AE_3_0[AE_3_0__T_530_addr]; // @[loaf.scala 147:67]
  assign AE_3_0__T_153_data = {slcBuf_e,slcBuf_a};
  assign AE_3_0__T_153_addr = prev_idx;
  assign AE_3_0__T_153_mask = 1'h1;
  assign AE_3_0__T_153_en = _T_2 ? _GEN_1109 : 1'h0;
  assign AE_3_1__T_618_addr = _T_494 + _GEN_4796;
  assign AE_3_1__T_618_data = AE_3_1[AE_3_1__T_618_addr]; // @[loaf.scala 147:67]
  assign AE_3_1__T_159_data = {slcBuf_e,slcBuf_a};
  assign AE_3_1__T_159_addr = prev_idx;
  assign AE_3_1__T_159_mask = 1'h1;
  assign AE_3_1__T_159_en = _T_2 ? _GEN_1114 : 1'h0;
  assign AE_3_2__T_706_addr = _T_494 + _GEN_4796;
  assign AE_3_2__T_706_data = AE_3_2[AE_3_2__T_706_addr]; // @[loaf.scala 147:67]
  assign AE_3_2__T_165_data = {slcBuf_e,slcBuf_a};
  assign AE_3_2__T_165_addr = prev_idx;
  assign AE_3_2__T_165_mask = 1'h1;
  assign AE_3_2__T_165_en = _T_2 ? _GEN_1119 : 1'h0;
  assign AE_3_3__T_794_addr = _T_494 + _GEN_4796;
  assign AE_3_3__T_794_data = AE_3_3[AE_3_3__T_794_addr]; // @[loaf.scala 147:67]
  assign AE_3_3__T_171_data = {slcBuf_e,slcBuf_a};
  assign AE_3_3__T_171_addr = prev_idx;
  assign AE_3_3__T_171_mask = 1'h1;
  assign AE_3_3__T_171_en = _T_2 ? _GEN_1124 : 1'h0;
  assign AE_3_4__T_882_addr = _T_494 + _GEN_4796;
  assign AE_3_4__T_882_data = AE_3_4[AE_3_4__T_882_addr]; // @[loaf.scala 147:67]
  assign AE_3_4__T_177_data = {slcBuf_e,slcBuf_a};
  assign AE_3_4__T_177_addr = prev_idx;
  assign AE_3_4__T_177_mask = 1'h1;
  assign AE_3_4__T_177_en = _T_2 ? _GEN_1129 : 1'h0;
  assign AE_3_5__T_970_addr = _T_494 + _GEN_4796;
  assign AE_3_5__T_970_data = AE_3_5[AE_3_5__T_970_addr]; // @[loaf.scala 147:67]
  assign AE_3_5__T_183_data = {slcBuf_e,slcBuf_a};
  assign AE_3_5__T_183_addr = prev_idx;
  assign AE_3_5__T_183_mask = 1'h1;
  assign AE_3_5__T_183_en = _T_2 ? _GEN_1134 : 1'h0;
  assign AE_3_6__T_1058_addr = _T_494 + _GEN_4796;
  assign AE_3_6__T_1058_data = AE_3_6[AE_3_6__T_1058_addr]; // @[loaf.scala 147:67]
  assign AE_3_6__T_189_data = {slcBuf_e,slcBuf_a};
  assign AE_3_6__T_189_addr = prev_idx;
  assign AE_3_6__T_189_mask = 1'h1;
  assign AE_3_6__T_189_en = _T_2 ? _GEN_1139 : 1'h0;
  assign AE_3_7__T_1146_addr = _T_494 + _GEN_4796;
  assign AE_3_7__T_1146_data = AE_3_7[AE_3_7__T_1146_addr]; // @[loaf.scala 147:67]
  assign AE_3_7__T_195_data = {slcBuf_e,slcBuf_a};
  assign AE_3_7__T_195_addr = prev_idx;
  assign AE_3_7__T_195_mask = 1'h1;
  assign AE_3_7__T_195_en = _T_2 ? _GEN_1144 : 1'h0;
  assign AE_4_0__T_541_addr = _T_494 + _GEN_4796;
  assign AE_4_0__T_541_data = AE_4_0[AE_4_0__T_541_addr]; // @[loaf.scala 147:67]
  assign AE_4_0__T_201_data = {slcBuf_e,slcBuf_a};
  assign AE_4_0__T_201_addr = prev_idx;
  assign AE_4_0__T_201_mask = 1'h1;
  assign AE_4_0__T_201_en = _T_2 ? _GEN_1149 : 1'h0;
  assign AE_4_1__T_629_addr = _T_494 + _GEN_4796;
  assign AE_4_1__T_629_data = AE_4_1[AE_4_1__T_629_addr]; // @[loaf.scala 147:67]
  assign AE_4_1__T_207_data = {slcBuf_e,slcBuf_a};
  assign AE_4_1__T_207_addr = prev_idx;
  assign AE_4_1__T_207_mask = 1'h1;
  assign AE_4_1__T_207_en = _T_2 ? _GEN_1154 : 1'h0;
  assign AE_4_2__T_717_addr = _T_494 + _GEN_4796;
  assign AE_4_2__T_717_data = AE_4_2[AE_4_2__T_717_addr]; // @[loaf.scala 147:67]
  assign AE_4_2__T_213_data = {slcBuf_e,slcBuf_a};
  assign AE_4_2__T_213_addr = prev_idx;
  assign AE_4_2__T_213_mask = 1'h1;
  assign AE_4_2__T_213_en = _T_2 ? _GEN_1159 : 1'h0;
  assign AE_4_3__T_805_addr = _T_494 + _GEN_4796;
  assign AE_4_3__T_805_data = AE_4_3[AE_4_3__T_805_addr]; // @[loaf.scala 147:67]
  assign AE_4_3__T_219_data = {slcBuf_e,slcBuf_a};
  assign AE_4_3__T_219_addr = prev_idx;
  assign AE_4_3__T_219_mask = 1'h1;
  assign AE_4_3__T_219_en = _T_2 ? _GEN_1164 : 1'h0;
  assign AE_4_4__T_893_addr = _T_494 + _GEN_4796;
  assign AE_4_4__T_893_data = AE_4_4[AE_4_4__T_893_addr]; // @[loaf.scala 147:67]
  assign AE_4_4__T_225_data = {slcBuf_e,slcBuf_a};
  assign AE_4_4__T_225_addr = prev_idx;
  assign AE_4_4__T_225_mask = 1'h1;
  assign AE_4_4__T_225_en = _T_2 ? _GEN_1169 : 1'h0;
  assign AE_4_5__T_981_addr = _T_494 + _GEN_4796;
  assign AE_4_5__T_981_data = AE_4_5[AE_4_5__T_981_addr]; // @[loaf.scala 147:67]
  assign AE_4_5__T_231_data = {slcBuf_e,slcBuf_a};
  assign AE_4_5__T_231_addr = prev_idx;
  assign AE_4_5__T_231_mask = 1'h1;
  assign AE_4_5__T_231_en = _T_2 ? _GEN_1174 : 1'h0;
  assign AE_4_6__T_1069_addr = _T_494 + _GEN_4796;
  assign AE_4_6__T_1069_data = AE_4_6[AE_4_6__T_1069_addr]; // @[loaf.scala 147:67]
  assign AE_4_6__T_237_data = {slcBuf_e,slcBuf_a};
  assign AE_4_6__T_237_addr = prev_idx;
  assign AE_4_6__T_237_mask = 1'h1;
  assign AE_4_6__T_237_en = _T_2 ? _GEN_1179 : 1'h0;
  assign AE_4_7__T_1157_addr = _T_494 + _GEN_4796;
  assign AE_4_7__T_1157_data = AE_4_7[AE_4_7__T_1157_addr]; // @[loaf.scala 147:67]
  assign AE_4_7__T_243_data = {slcBuf_e,slcBuf_a};
  assign AE_4_7__T_243_addr = prev_idx;
  assign AE_4_7__T_243_mask = 1'h1;
  assign AE_4_7__T_243_en = _T_2 ? _GEN_1184 : 1'h0;
  assign AE_5_0__T_552_addr = _T_494 + _GEN_4796;
  assign AE_5_0__T_552_data = AE_5_0[AE_5_0__T_552_addr]; // @[loaf.scala 147:67]
  assign AE_5_0__T_249_data = {slcBuf_e,slcBuf_a};
  assign AE_5_0__T_249_addr = prev_idx;
  assign AE_5_0__T_249_mask = 1'h1;
  assign AE_5_0__T_249_en = _T_2 ? _GEN_1189 : 1'h0;
  assign AE_5_1__T_640_addr = _T_494 + _GEN_4796;
  assign AE_5_1__T_640_data = AE_5_1[AE_5_1__T_640_addr]; // @[loaf.scala 147:67]
  assign AE_5_1__T_255_data = {slcBuf_e,slcBuf_a};
  assign AE_5_1__T_255_addr = prev_idx;
  assign AE_5_1__T_255_mask = 1'h1;
  assign AE_5_1__T_255_en = _T_2 ? _GEN_1194 : 1'h0;
  assign AE_5_2__T_728_addr = _T_494 + _GEN_4796;
  assign AE_5_2__T_728_data = AE_5_2[AE_5_2__T_728_addr]; // @[loaf.scala 147:67]
  assign AE_5_2__T_261_data = {slcBuf_e,slcBuf_a};
  assign AE_5_2__T_261_addr = prev_idx;
  assign AE_5_2__T_261_mask = 1'h1;
  assign AE_5_2__T_261_en = _T_2 ? _GEN_1199 : 1'h0;
  assign AE_5_3__T_816_addr = _T_494 + _GEN_4796;
  assign AE_5_3__T_816_data = AE_5_3[AE_5_3__T_816_addr]; // @[loaf.scala 147:67]
  assign AE_5_3__T_267_data = {slcBuf_e,slcBuf_a};
  assign AE_5_3__T_267_addr = prev_idx;
  assign AE_5_3__T_267_mask = 1'h1;
  assign AE_5_3__T_267_en = _T_2 ? _GEN_1204 : 1'h0;
  assign AE_5_4__T_904_addr = _T_494 + _GEN_4796;
  assign AE_5_4__T_904_data = AE_5_4[AE_5_4__T_904_addr]; // @[loaf.scala 147:67]
  assign AE_5_4__T_273_data = {slcBuf_e,slcBuf_a};
  assign AE_5_4__T_273_addr = prev_idx;
  assign AE_5_4__T_273_mask = 1'h1;
  assign AE_5_4__T_273_en = _T_2 ? _GEN_1209 : 1'h0;
  assign AE_5_5__T_992_addr = _T_494 + _GEN_4796;
  assign AE_5_5__T_992_data = AE_5_5[AE_5_5__T_992_addr]; // @[loaf.scala 147:67]
  assign AE_5_5__T_279_data = {slcBuf_e,slcBuf_a};
  assign AE_5_5__T_279_addr = prev_idx;
  assign AE_5_5__T_279_mask = 1'h1;
  assign AE_5_5__T_279_en = _T_2 ? _GEN_1214 : 1'h0;
  assign AE_5_6__T_1080_addr = _T_494 + _GEN_4796;
  assign AE_5_6__T_1080_data = AE_5_6[AE_5_6__T_1080_addr]; // @[loaf.scala 147:67]
  assign AE_5_6__T_285_data = {slcBuf_e,slcBuf_a};
  assign AE_5_6__T_285_addr = prev_idx;
  assign AE_5_6__T_285_mask = 1'h1;
  assign AE_5_6__T_285_en = _T_2 ? _GEN_1219 : 1'h0;
  assign AE_5_7__T_1168_addr = _T_494 + _GEN_4796;
  assign AE_5_7__T_1168_data = AE_5_7[AE_5_7__T_1168_addr]; // @[loaf.scala 147:67]
  assign AE_5_7__T_291_data = {slcBuf_e,slcBuf_a};
  assign AE_5_7__T_291_addr = prev_idx;
  assign AE_5_7__T_291_mask = 1'h1;
  assign AE_5_7__T_291_en = _T_2 ? _GEN_1224 : 1'h0;
  assign AE_6_0__T_563_addr = _T_494 + _GEN_4796;
  assign AE_6_0__T_563_data = AE_6_0[AE_6_0__T_563_addr]; // @[loaf.scala 147:67]
  assign AE_6_0__T_297_data = {slcBuf_e,slcBuf_a};
  assign AE_6_0__T_297_addr = prev_idx;
  assign AE_6_0__T_297_mask = 1'h1;
  assign AE_6_0__T_297_en = _T_2 ? _GEN_1229 : 1'h0;
  assign AE_6_1__T_651_addr = _T_494 + _GEN_4796;
  assign AE_6_1__T_651_data = AE_6_1[AE_6_1__T_651_addr]; // @[loaf.scala 147:67]
  assign AE_6_1__T_303_data = {slcBuf_e,slcBuf_a};
  assign AE_6_1__T_303_addr = prev_idx;
  assign AE_6_1__T_303_mask = 1'h1;
  assign AE_6_1__T_303_en = _T_2 ? _GEN_1234 : 1'h0;
  assign AE_6_2__T_739_addr = _T_494 + _GEN_4796;
  assign AE_6_2__T_739_data = AE_6_2[AE_6_2__T_739_addr]; // @[loaf.scala 147:67]
  assign AE_6_2__T_309_data = {slcBuf_e,slcBuf_a};
  assign AE_6_2__T_309_addr = prev_idx;
  assign AE_6_2__T_309_mask = 1'h1;
  assign AE_6_2__T_309_en = _T_2 ? _GEN_1239 : 1'h0;
  assign AE_6_3__T_827_addr = _T_494 + _GEN_4796;
  assign AE_6_3__T_827_data = AE_6_3[AE_6_3__T_827_addr]; // @[loaf.scala 147:67]
  assign AE_6_3__T_315_data = {slcBuf_e,slcBuf_a};
  assign AE_6_3__T_315_addr = prev_idx;
  assign AE_6_3__T_315_mask = 1'h1;
  assign AE_6_3__T_315_en = _T_2 ? _GEN_1244 : 1'h0;
  assign AE_6_4__T_915_addr = _T_494 + _GEN_4796;
  assign AE_6_4__T_915_data = AE_6_4[AE_6_4__T_915_addr]; // @[loaf.scala 147:67]
  assign AE_6_4__T_321_data = {slcBuf_e,slcBuf_a};
  assign AE_6_4__T_321_addr = prev_idx;
  assign AE_6_4__T_321_mask = 1'h1;
  assign AE_6_4__T_321_en = _T_2 ? _GEN_1249 : 1'h0;
  assign AE_6_5__T_1003_addr = _T_494 + _GEN_4796;
  assign AE_6_5__T_1003_data = AE_6_5[AE_6_5__T_1003_addr]; // @[loaf.scala 147:67]
  assign AE_6_5__T_327_data = {slcBuf_e,slcBuf_a};
  assign AE_6_5__T_327_addr = prev_idx;
  assign AE_6_5__T_327_mask = 1'h1;
  assign AE_6_5__T_327_en = _T_2 ? _GEN_1254 : 1'h0;
  assign AE_6_6__T_1091_addr = _T_494 + _GEN_4796;
  assign AE_6_6__T_1091_data = AE_6_6[AE_6_6__T_1091_addr]; // @[loaf.scala 147:67]
  assign AE_6_6__T_333_data = {slcBuf_e,slcBuf_a};
  assign AE_6_6__T_333_addr = prev_idx;
  assign AE_6_6__T_333_mask = 1'h1;
  assign AE_6_6__T_333_en = _T_2 ? _GEN_1259 : 1'h0;
  assign AE_6_7__T_1179_addr = _T_494 + _GEN_4796;
  assign AE_6_7__T_1179_data = AE_6_7[AE_6_7__T_1179_addr]; // @[loaf.scala 147:67]
  assign AE_6_7__T_339_data = {slcBuf_e,slcBuf_a};
  assign AE_6_7__T_339_addr = prev_idx;
  assign AE_6_7__T_339_mask = 1'h1;
  assign AE_6_7__T_339_en = _T_2 ? _GEN_1264 : 1'h0;
  assign AE_7_0__T_574_addr = _T_494 + _GEN_4796;
  assign AE_7_0__T_574_data = AE_7_0[AE_7_0__T_574_addr]; // @[loaf.scala 147:67]
  assign AE_7_0__T_345_data = {slcBuf_e,slcBuf_a};
  assign AE_7_0__T_345_addr = prev_idx;
  assign AE_7_0__T_345_mask = 1'h1;
  assign AE_7_0__T_345_en = _T_2 ? _GEN_1269 : 1'h0;
  assign AE_7_1__T_662_addr = _T_494 + _GEN_4796;
  assign AE_7_1__T_662_data = AE_7_1[AE_7_1__T_662_addr]; // @[loaf.scala 147:67]
  assign AE_7_1__T_351_data = {slcBuf_e,slcBuf_a};
  assign AE_7_1__T_351_addr = prev_idx;
  assign AE_7_1__T_351_mask = 1'h1;
  assign AE_7_1__T_351_en = _T_2 ? _GEN_1274 : 1'h0;
  assign AE_7_2__T_750_addr = _T_494 + _GEN_4796;
  assign AE_7_2__T_750_data = AE_7_2[AE_7_2__T_750_addr]; // @[loaf.scala 147:67]
  assign AE_7_2__T_357_data = {slcBuf_e,slcBuf_a};
  assign AE_7_2__T_357_addr = prev_idx;
  assign AE_7_2__T_357_mask = 1'h1;
  assign AE_7_2__T_357_en = _T_2 ? _GEN_1279 : 1'h0;
  assign AE_7_3__T_838_addr = _T_494 + _GEN_4796;
  assign AE_7_3__T_838_data = AE_7_3[AE_7_3__T_838_addr]; // @[loaf.scala 147:67]
  assign AE_7_3__T_363_data = {slcBuf_e,slcBuf_a};
  assign AE_7_3__T_363_addr = prev_idx;
  assign AE_7_3__T_363_mask = 1'h1;
  assign AE_7_3__T_363_en = _T_2 ? _GEN_1284 : 1'h0;
  assign AE_7_4__T_926_addr = _T_494 + _GEN_4796;
  assign AE_7_4__T_926_data = AE_7_4[AE_7_4__T_926_addr]; // @[loaf.scala 147:67]
  assign AE_7_4__T_369_data = {slcBuf_e,slcBuf_a};
  assign AE_7_4__T_369_addr = prev_idx;
  assign AE_7_4__T_369_mask = 1'h1;
  assign AE_7_4__T_369_en = _T_2 ? _GEN_1289 : 1'h0;
  assign AE_7_5__T_1014_addr = _T_494 + _GEN_4796;
  assign AE_7_5__T_1014_data = AE_7_5[AE_7_5__T_1014_addr]; // @[loaf.scala 147:67]
  assign AE_7_5__T_375_data = {slcBuf_e,slcBuf_a};
  assign AE_7_5__T_375_addr = prev_idx;
  assign AE_7_5__T_375_mask = 1'h1;
  assign AE_7_5__T_375_en = _T_2 ? _GEN_1294 : 1'h0;
  assign AE_7_6__T_1102_addr = _T_494 + _GEN_4796;
  assign AE_7_6__T_1102_data = AE_7_6[AE_7_6__T_1102_addr]; // @[loaf.scala 147:67]
  assign AE_7_6__T_381_data = {slcBuf_e,slcBuf_a};
  assign AE_7_6__T_381_addr = prev_idx;
  assign AE_7_6__T_381_mask = 1'h1;
  assign AE_7_6__T_381_en = _T_2 ? _GEN_1299 : 1'h0;
  assign AE_7_7__T_1190_addr = _T_494 + _GEN_4796;
  assign AE_7_7__T_1190_data = AE_7_7[AE_7_7__T_1190_addr]; // @[loaf.scala 147:67]
  assign AE_7_7__T_387_data = {slcBuf_e,slcBuf_a};
  assign AE_7_7__T_387_addr = prev_idx;
  assign AE_7_7__T_387_mask = 1'h1;
  assign AE_7_7__T_387_en = _T_2 ? _GEN_1304 : 1'h0;
  assign _T_1 = doneLoading == 1'h0; // @[loaf.scala 170:22]
  assign _T_2 = io_start & _T_1; // @[loaf.scala 170:19]
  assign _T_3 = io_slc_valid | lastLoad; // @[loaf.scala 174:27]
  assign _T_4 = 3'h0 == prev_lo_i; // @[loaf.scala 179:24]
  assign _T_5 = 3'h0 == prev_lo_j; // @[loaf.scala 179:45]
  assign _T_6 = _T_4 & _T_5; // @[loaf.scala 179:38]
  assign _T_11 = 3'h1 == prev_lo_j; // @[loaf.scala 179:45]
  assign _T_12 = _T_4 & _T_11; // @[loaf.scala 179:38]
  assign _T_17 = 3'h2 == prev_lo_j; // @[loaf.scala 179:45]
  assign _T_18 = _T_4 & _T_17; // @[loaf.scala 179:38]
  assign _T_23 = 3'h3 == prev_lo_j; // @[loaf.scala 179:45]
  assign _T_24 = _T_4 & _T_23; // @[loaf.scala 179:38]
  assign _T_29 = 3'h4 == prev_lo_j; // @[loaf.scala 179:45]
  assign _T_30 = _T_4 & _T_29; // @[loaf.scala 179:38]
  assign _T_35 = 3'h5 == prev_lo_j; // @[loaf.scala 179:45]
  assign _T_36 = _T_4 & _T_35; // @[loaf.scala 179:38]
  assign _T_41 = 3'h6 == prev_lo_j; // @[loaf.scala 179:45]
  assign _T_42 = _T_4 & _T_41; // @[loaf.scala 179:38]
  assign _T_47 = 3'h7 == prev_lo_j; // @[loaf.scala 179:45]
  assign _T_48 = _T_4 & _T_47; // @[loaf.scala 179:38]
  assign _T_52 = 3'h1 == prev_lo_i; // @[loaf.scala 179:24]
  assign _T_54 = _T_52 & _T_5; // @[loaf.scala 179:38]
  assign _T_60 = _T_52 & _T_11; // @[loaf.scala 179:38]
  assign _T_66 = _T_52 & _T_17; // @[loaf.scala 179:38]
  assign _T_72 = _T_52 & _T_23; // @[loaf.scala 179:38]
  assign _T_78 = _T_52 & _T_29; // @[loaf.scala 179:38]
  assign _T_84 = _T_52 & _T_35; // @[loaf.scala 179:38]
  assign _T_90 = _T_52 & _T_41; // @[loaf.scala 179:38]
  assign _T_96 = _T_52 & _T_47; // @[loaf.scala 179:38]
  assign _T_100 = 3'h2 == prev_lo_i; // @[loaf.scala 179:24]
  assign _T_102 = _T_100 & _T_5; // @[loaf.scala 179:38]
  assign _T_108 = _T_100 & _T_11; // @[loaf.scala 179:38]
  assign _T_114 = _T_100 & _T_17; // @[loaf.scala 179:38]
  assign _T_120 = _T_100 & _T_23; // @[loaf.scala 179:38]
  assign _T_126 = _T_100 & _T_29; // @[loaf.scala 179:38]
  assign _T_132 = _T_100 & _T_35; // @[loaf.scala 179:38]
  assign _T_138 = _T_100 & _T_41; // @[loaf.scala 179:38]
  assign _T_144 = _T_100 & _T_47; // @[loaf.scala 179:38]
  assign _T_148 = 3'h3 == prev_lo_i; // @[loaf.scala 179:24]
  assign _T_150 = _T_148 & _T_5; // @[loaf.scala 179:38]
  assign _T_156 = _T_148 & _T_11; // @[loaf.scala 179:38]
  assign _T_162 = _T_148 & _T_17; // @[loaf.scala 179:38]
  assign _T_168 = _T_148 & _T_23; // @[loaf.scala 179:38]
  assign _T_174 = _T_148 & _T_29; // @[loaf.scala 179:38]
  assign _T_180 = _T_148 & _T_35; // @[loaf.scala 179:38]
  assign _T_186 = _T_148 & _T_41; // @[loaf.scala 179:38]
  assign _T_192 = _T_148 & _T_47; // @[loaf.scala 179:38]
  assign _T_196 = 3'h4 == prev_lo_i; // @[loaf.scala 179:24]
  assign _T_198 = _T_196 & _T_5; // @[loaf.scala 179:38]
  assign _T_204 = _T_196 & _T_11; // @[loaf.scala 179:38]
  assign _T_210 = _T_196 & _T_17; // @[loaf.scala 179:38]
  assign _T_216 = _T_196 & _T_23; // @[loaf.scala 179:38]
  assign _T_222 = _T_196 & _T_29; // @[loaf.scala 179:38]
  assign _T_228 = _T_196 & _T_35; // @[loaf.scala 179:38]
  assign _T_234 = _T_196 & _T_41; // @[loaf.scala 179:38]
  assign _T_240 = _T_196 & _T_47; // @[loaf.scala 179:38]
  assign _T_244 = 3'h5 == prev_lo_i; // @[loaf.scala 179:24]
  assign _T_246 = _T_244 & _T_5; // @[loaf.scala 179:38]
  assign _T_252 = _T_244 & _T_11; // @[loaf.scala 179:38]
  assign _T_258 = _T_244 & _T_17; // @[loaf.scala 179:38]
  assign _T_264 = _T_244 & _T_23; // @[loaf.scala 179:38]
  assign _T_270 = _T_244 & _T_29; // @[loaf.scala 179:38]
  assign _T_276 = _T_244 & _T_35; // @[loaf.scala 179:38]
  assign _T_282 = _T_244 & _T_41; // @[loaf.scala 179:38]
  assign _T_288 = _T_244 & _T_47; // @[loaf.scala 179:38]
  assign _T_292 = 3'h6 == prev_lo_i; // @[loaf.scala 179:24]
  assign _T_294 = _T_292 & _T_5; // @[loaf.scala 179:38]
  assign _T_300 = _T_292 & _T_11; // @[loaf.scala 179:38]
  assign _T_306 = _T_292 & _T_17; // @[loaf.scala 179:38]
  assign _T_312 = _T_292 & _T_23; // @[loaf.scala 179:38]
  assign _T_318 = _T_292 & _T_29; // @[loaf.scala 179:38]
  assign _T_324 = _T_292 & _T_35; // @[loaf.scala 179:38]
  assign _T_330 = _T_292 & _T_41; // @[loaf.scala 179:38]
  assign _T_336 = _T_292 & _T_47; // @[loaf.scala 179:38]
  assign _T_340 = 3'h7 == prev_lo_i; // @[loaf.scala 179:24]
  assign _T_342 = _T_340 & _T_5; // @[loaf.scala 179:38]
  assign _T_348 = _T_340 & _T_11; // @[loaf.scala 179:38]
  assign _T_354 = _T_340 & _T_17; // @[loaf.scala 179:38]
  assign _T_360 = _T_340 & _T_23; // @[loaf.scala 179:38]
  assign _T_366 = _T_340 & _T_29; // @[loaf.scala 179:38]
  assign _T_372 = _T_340 & _T_35; // @[loaf.scala 179:38]
  assign _T_378 = _T_340 & _T_41; // @[loaf.scala 179:38]
  assign _T_384 = _T_340 & _T_47; // @[loaf.scala 179:38]
  assign _GEN_322 = slcValid ? _T_6 : 1'h0; // @[loaf.scala 176:26]
  assign _GEN_327 = slcValid ? _T_12 : 1'h0; // @[loaf.scala 176:26]
  assign _GEN_332 = slcValid ? _T_18 : 1'h0; // @[loaf.scala 176:26]
  assign _GEN_337 = slcValid ? _T_24 : 1'h0; // @[loaf.scala 176:26]
  assign _GEN_342 = slcValid ? _T_30 : 1'h0; // @[loaf.scala 176:26]
  assign _GEN_347 = slcValid ? _T_36 : 1'h0; // @[loaf.scala 176:26]
  assign _GEN_352 = slcValid ? _T_42 : 1'h0; // @[loaf.scala 176:26]
  assign _GEN_357 = slcValid ? _T_48 : 1'h0; // @[loaf.scala 176:26]
  assign _GEN_362 = slcValid ? _T_54 : 1'h0; // @[loaf.scala 176:26]
  assign _GEN_367 = slcValid ? _T_60 : 1'h0; // @[loaf.scala 176:26]
  assign _GEN_372 = slcValid ? _T_66 : 1'h0; // @[loaf.scala 176:26]
  assign _GEN_377 = slcValid ? _T_72 : 1'h0; // @[loaf.scala 176:26]
  assign _GEN_382 = slcValid ? _T_78 : 1'h0; // @[loaf.scala 176:26]
  assign _GEN_387 = slcValid ? _T_84 : 1'h0; // @[loaf.scala 176:26]
  assign _GEN_392 = slcValid ? _T_90 : 1'h0; // @[loaf.scala 176:26]
  assign _GEN_397 = slcValid ? _T_96 : 1'h0; // @[loaf.scala 176:26]
  assign _GEN_402 = slcValid ? _T_102 : 1'h0; // @[loaf.scala 176:26]
  assign _GEN_407 = slcValid ? _T_108 : 1'h0; // @[loaf.scala 176:26]
  assign _GEN_412 = slcValid ? _T_114 : 1'h0; // @[loaf.scala 176:26]
  assign _GEN_417 = slcValid ? _T_120 : 1'h0; // @[loaf.scala 176:26]
  assign _GEN_422 = slcValid ? _T_126 : 1'h0; // @[loaf.scala 176:26]
  assign _GEN_427 = slcValid ? _T_132 : 1'h0; // @[loaf.scala 176:26]
  assign _GEN_432 = slcValid ? _T_138 : 1'h0; // @[loaf.scala 176:26]
  assign _GEN_437 = slcValid ? _T_144 : 1'h0; // @[loaf.scala 176:26]
  assign _GEN_442 = slcValid ? _T_150 : 1'h0; // @[loaf.scala 176:26]
  assign _GEN_447 = slcValid ? _T_156 : 1'h0; // @[loaf.scala 176:26]
  assign _GEN_452 = slcValid ? _T_162 : 1'h0; // @[loaf.scala 176:26]
  assign _GEN_457 = slcValid ? _T_168 : 1'h0; // @[loaf.scala 176:26]
  assign _GEN_462 = slcValid ? _T_174 : 1'h0; // @[loaf.scala 176:26]
  assign _GEN_467 = slcValid ? _T_180 : 1'h0; // @[loaf.scala 176:26]
  assign _GEN_472 = slcValid ? _T_186 : 1'h0; // @[loaf.scala 176:26]
  assign _GEN_477 = slcValid ? _T_192 : 1'h0; // @[loaf.scala 176:26]
  assign _GEN_482 = slcValid ? _T_198 : 1'h0; // @[loaf.scala 176:26]
  assign _GEN_487 = slcValid ? _T_204 : 1'h0; // @[loaf.scala 176:26]
  assign _GEN_492 = slcValid ? _T_210 : 1'h0; // @[loaf.scala 176:26]
  assign _GEN_497 = slcValid ? _T_216 : 1'h0; // @[loaf.scala 176:26]
  assign _GEN_502 = slcValid ? _T_222 : 1'h0; // @[loaf.scala 176:26]
  assign _GEN_507 = slcValid ? _T_228 : 1'h0; // @[loaf.scala 176:26]
  assign _GEN_512 = slcValid ? _T_234 : 1'h0; // @[loaf.scala 176:26]
  assign _GEN_517 = slcValid ? _T_240 : 1'h0; // @[loaf.scala 176:26]
  assign _GEN_522 = slcValid ? _T_246 : 1'h0; // @[loaf.scala 176:26]
  assign _GEN_527 = slcValid ? _T_252 : 1'h0; // @[loaf.scala 176:26]
  assign _GEN_532 = slcValid ? _T_258 : 1'h0; // @[loaf.scala 176:26]
  assign _GEN_537 = slcValid ? _T_264 : 1'h0; // @[loaf.scala 176:26]
  assign _GEN_542 = slcValid ? _T_270 : 1'h0; // @[loaf.scala 176:26]
  assign _GEN_547 = slcValid ? _T_276 : 1'h0; // @[loaf.scala 176:26]
  assign _GEN_552 = slcValid ? _T_282 : 1'h0; // @[loaf.scala 176:26]
  assign _GEN_557 = slcValid ? _T_288 : 1'h0; // @[loaf.scala 176:26]
  assign _GEN_562 = slcValid ? _T_294 : 1'h0; // @[loaf.scala 176:26]
  assign _GEN_567 = slcValid ? _T_300 : 1'h0; // @[loaf.scala 176:26]
  assign _GEN_572 = slcValid ? _T_306 : 1'h0; // @[loaf.scala 176:26]
  assign _GEN_577 = slcValid ? _T_312 : 1'h0; // @[loaf.scala 176:26]
  assign _GEN_582 = slcValid ? _T_318 : 1'h0; // @[loaf.scala 176:26]
  assign _GEN_587 = slcValid ? _T_324 : 1'h0; // @[loaf.scala 176:26]
  assign _GEN_592 = slcValid ? _T_330 : 1'h0; // @[loaf.scala 176:26]
  assign _GEN_597 = slcValid ? _T_336 : 1'h0; // @[loaf.scala 176:26]
  assign _GEN_602 = slcValid ? _T_342 : 1'h0; // @[loaf.scala 176:26]
  assign _GEN_607 = slcValid ? _T_348 : 1'h0; // @[loaf.scala 176:26]
  assign _GEN_612 = slcValid ? _T_354 : 1'h0; // @[loaf.scala 176:26]
  assign _GEN_617 = slcValid ? _T_360 : 1'h0; // @[loaf.scala 176:26]
  assign _GEN_622 = slcValid ? _T_366 : 1'h0; // @[loaf.scala 176:26]
  assign _GEN_627 = slcValid ? _T_372 : 1'h0; // @[loaf.scala 176:26]
  assign _GEN_632 = slcValid ? _T_378 : 1'h0; // @[loaf.scala 176:26]
  assign _GEN_637 = slcValid ? _T_384 : 1'h0; // @[loaf.scala 176:26]
  assign _T_388 = load_i[2:0]; // @[loaf.scala 193:19]
  assign _T_389 = load_i[4:3]; // @[loaf.scala 195:28]
  assign _T_390 = load_j[2:0]; // @[loaf.scala 197:19]
  assign _T_391 = load_j[4:3]; // @[loaf.scala 199:28]
  assign _T_392 = {io_loadIdx, 4'h0}; // @[loaf.scala 201:32]
  assign _T_393 = {_T_389, 2'h0}; // @[loaf.scala 201:68]
  assign _GEN_4793 = {{1'd0}, _T_393}; // @[loaf.scala 201:59]
  assign _T_395 = _T_392 + _GEN_4793; // @[loaf.scala 201:59]
  assign _GEN_4794 = {{3'd0}, _T_391}; // @[loaf.scala 201:92]
  assign _T_397 = _T_395 + _GEN_4794; // @[loaf.scala 201:92]
  assign _T_398 = load_j != 5'h17; // @[loaf.scala 209:25]
  assign _T_400 = load_j + 5'h1; // @[loaf.scala 210:30]
  assign _T_401 = load_i != 5'h17; // @[loaf.scala 213:27]
  assign _T_403 = load_i + 5'h1; // @[loaf.scala 214:32]
  assign _GEN_647 = lastLoad ? 1'h0 : 1'h1; // @[loaf.scala 185:26]
  assign _GEN_658 = _T_3 ? _GEN_322 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_663 = _T_3 ? _GEN_327 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_668 = _T_3 ? _GEN_332 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_673 = _T_3 ? _GEN_337 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_678 = _T_3 ? _GEN_342 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_683 = _T_3 ? _GEN_347 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_688 = _T_3 ? _GEN_352 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_693 = _T_3 ? _GEN_357 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_698 = _T_3 ? _GEN_362 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_703 = _T_3 ? _GEN_367 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_708 = _T_3 ? _GEN_372 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_713 = _T_3 ? _GEN_377 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_718 = _T_3 ? _GEN_382 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_723 = _T_3 ? _GEN_387 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_728 = _T_3 ? _GEN_392 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_733 = _T_3 ? _GEN_397 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_738 = _T_3 ? _GEN_402 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_743 = _T_3 ? _GEN_407 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_748 = _T_3 ? _GEN_412 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_753 = _T_3 ? _GEN_417 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_758 = _T_3 ? _GEN_422 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_763 = _T_3 ? _GEN_427 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_768 = _T_3 ? _GEN_432 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_773 = _T_3 ? _GEN_437 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_778 = _T_3 ? _GEN_442 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_783 = _T_3 ? _GEN_447 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_788 = _T_3 ? _GEN_452 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_793 = _T_3 ? _GEN_457 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_798 = _T_3 ? _GEN_462 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_803 = _T_3 ? _GEN_467 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_808 = _T_3 ? _GEN_472 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_813 = _T_3 ? _GEN_477 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_818 = _T_3 ? _GEN_482 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_823 = _T_3 ? _GEN_487 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_828 = _T_3 ? _GEN_492 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_833 = _T_3 ? _GEN_497 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_838 = _T_3 ? _GEN_502 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_843 = _T_3 ? _GEN_507 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_848 = _T_3 ? _GEN_512 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_853 = _T_3 ? _GEN_517 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_858 = _T_3 ? _GEN_522 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_863 = _T_3 ? _GEN_527 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_868 = _T_3 ? _GEN_532 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_873 = _T_3 ? _GEN_537 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_878 = _T_3 ? _GEN_542 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_883 = _T_3 ? _GEN_547 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_888 = _T_3 ? _GEN_552 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_893 = _T_3 ? _GEN_557 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_898 = _T_3 ? _GEN_562 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_903 = _T_3 ? _GEN_567 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_908 = _T_3 ? _GEN_572 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_913 = _T_3 ? _GEN_577 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_918 = _T_3 ? _GEN_582 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_923 = _T_3 ? _GEN_587 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_928 = _T_3 ? _GEN_592 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_933 = _T_3 ? _GEN_597 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_938 = _T_3 ? _GEN_602 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_943 = _T_3 ? _GEN_607 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_948 = _T_3 ? _GEN_612 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_953 = _T_3 ? _GEN_617 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_958 = _T_3 ? _GEN_622 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_963 = _T_3 ? _GEN_627 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_968 = _T_3 ? _GEN_632 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_973 = _T_3 ? _GEN_637 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_978 = _T_3 ? _GEN_647 : 1'h0; // @[loaf.scala 174:40]
  assign _GEN_989 = io_modeLoad ? _GEN_658 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_994 = io_modeLoad ? _GEN_663 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_999 = io_modeLoad ? _GEN_668 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_1004 = io_modeLoad ? _GEN_673 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_1009 = io_modeLoad ? _GEN_678 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_1014 = io_modeLoad ? _GEN_683 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_1019 = io_modeLoad ? _GEN_688 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_1024 = io_modeLoad ? _GEN_693 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_1029 = io_modeLoad ? _GEN_698 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_1034 = io_modeLoad ? _GEN_703 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_1039 = io_modeLoad ? _GEN_708 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_1044 = io_modeLoad ? _GEN_713 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_1049 = io_modeLoad ? _GEN_718 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_1054 = io_modeLoad ? _GEN_723 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_1059 = io_modeLoad ? _GEN_728 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_1064 = io_modeLoad ? _GEN_733 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_1069 = io_modeLoad ? _GEN_738 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_1074 = io_modeLoad ? _GEN_743 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_1079 = io_modeLoad ? _GEN_748 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_1084 = io_modeLoad ? _GEN_753 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_1089 = io_modeLoad ? _GEN_758 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_1094 = io_modeLoad ? _GEN_763 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_1099 = io_modeLoad ? _GEN_768 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_1104 = io_modeLoad ? _GEN_773 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_1109 = io_modeLoad ? _GEN_778 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_1114 = io_modeLoad ? _GEN_783 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_1119 = io_modeLoad ? _GEN_788 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_1124 = io_modeLoad ? _GEN_793 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_1129 = io_modeLoad ? _GEN_798 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_1134 = io_modeLoad ? _GEN_803 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_1139 = io_modeLoad ? _GEN_808 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_1144 = io_modeLoad ? _GEN_813 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_1149 = io_modeLoad ? _GEN_818 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_1154 = io_modeLoad ? _GEN_823 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_1159 = io_modeLoad ? _GEN_828 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_1164 = io_modeLoad ? _GEN_833 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_1169 = io_modeLoad ? _GEN_838 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_1174 = io_modeLoad ? _GEN_843 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_1179 = io_modeLoad ? _GEN_848 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_1184 = io_modeLoad ? _GEN_853 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_1189 = io_modeLoad ? _GEN_858 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_1194 = io_modeLoad ? _GEN_863 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_1199 = io_modeLoad ? _GEN_868 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_1204 = io_modeLoad ? _GEN_873 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_1209 = io_modeLoad ? _GEN_878 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_1214 = io_modeLoad ? _GEN_883 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_1219 = io_modeLoad ? _GEN_888 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_1224 = io_modeLoad ? _GEN_893 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_1229 = io_modeLoad ? _GEN_898 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_1234 = io_modeLoad ? _GEN_903 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_1239 = io_modeLoad ? _GEN_908 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_1244 = io_modeLoad ? _GEN_913 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_1249 = io_modeLoad ? _GEN_918 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_1254 = io_modeLoad ? _GEN_923 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_1259 = io_modeLoad ? _GEN_928 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_1264 = io_modeLoad ? _GEN_933 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_1269 = io_modeLoad ? _GEN_938 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_1274 = io_modeLoad ? _GEN_943 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_1279 = io_modeLoad ? _GEN_948 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_1284 = io_modeLoad ? _GEN_953 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_1289 = io_modeLoad ? _GEN_958 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_1294 = io_modeLoad ? _GEN_963 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_1299 = io_modeLoad ? _GEN_968 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_1304 = io_modeLoad ? _GEN_973 : 1'h0; // @[loaf.scala 172:25]
  assign _GEN_1309 = io_modeLoad ? _GEN_978 : 1'h0; // @[loaf.scala 172:25]
  assign _T_450 = done == 1'h0; // @[loaf.scala 234:22]
  assign _T_451 = io_start & _T_450; // @[loaf.scala 234:19]
  assign _T_452 = doneLoading & io_modeCompute; // @[loaf.scala 236:24]
  assign _T_453 = phase == 1'h0; // @[loaf.scala 244:34]
  assign _T_454 = c == 2'h0; // @[loaf.scala 244:47]
  assign _T_455 = _T_453 & _T_454; // @[loaf.scala 244:42]
  assign _T_456 = io_off_valid == 1'h0; // @[loaf.scala 244:59]
  assign _T_457 = r == 2'h0; // @[loaf.scala 244:79]
  assign _T_458 = io_lof_valid == 1'h0; // @[loaf.scala 244:90]
  assign _T_459 = _T_457 & _T_458; // @[loaf.scala 244:87]
  assign _T_460 = _T_456 | _T_459; // @[loaf.scala 244:73]
  assign _T_461 = _T_455 & _T_460; // @[loaf.scala 244:55]
  assign _T_462 = _T_434 == 1'h0; // @[loaf.scala 246:14]
  assign _T_463 = _T_462 | io_out_ready; // @[loaf.scala 246:32]
  assign _T_465 = _T_461 == 1'h0; // @[loaf.scala 248:46]
  assign _T_466 = _T_453 & _T_465; // @[loaf.scala 248:43]
  assign _T_468 = r == 2'h2; // @[loaf.scala 249:47]
  assign _T_469 = _T_453 & _T_468; // @[loaf.scala 249:42]
  assign _T_471 = _T_469 & _T_465; // @[loaf.scala 249:61]
  assign _T_474 = _T_453 & _T_457; // @[loaf.scala 250:43]
  assign _T_476 = _T_474 & _T_465; // @[loaf.scala 250:56]
  assign _GEN_1763 = _T_466 ? _T_454 : 1'h0; // @[loaf.scala 257:50]
  assign _T_485 = _T_455 & _T_457; // @[loaf.scala 267:43]
  assign _T_487 = _T_485 & _T_465; // @[loaf.scala 267:56]
  assign _T_491 = {io_computeIdx, 4'h0}; // @[loaf.scala 275:39]
  assign _T_492 = {r, 2'h0}; // @[loaf.scala 275:72]
  assign _GEN_4795 = {{1'd0}, _T_492}; // @[loaf.scala 275:66]
  assign _T_494 = _T_491 + _GEN_4795; // @[loaf.scala 275:66]
  assign _GEN_4796 = {{3'd0}, c}; // @[loaf.scala 275:96]
  assign _T_499 = AE_0_0__T_497_data;
  assign _T_500 = _T_499[15:0]; // @[loaf.scala 276:58]
  assign _T_501 = _T_499[31:16]; // @[loaf.scala 276:58]
  assign _T_510 = AE_1_0__T_508_data;
  assign _T_511 = _T_510[15:0]; // @[loaf.scala 276:58]
  assign _T_512 = _T_510[31:16]; // @[loaf.scala 276:58]
  assign _T_521 = AE_2_0__T_519_data;
  assign _T_522 = _T_521[15:0]; // @[loaf.scala 276:58]
  assign _T_523 = _T_521[31:16]; // @[loaf.scala 276:58]
  assign _T_532 = AE_3_0__T_530_data;
  assign _T_533 = _T_532[15:0]; // @[loaf.scala 276:58]
  assign _T_534 = _T_532[31:16]; // @[loaf.scala 276:58]
  assign _T_543 = AE_4_0__T_541_data;
  assign _T_544 = _T_543[15:0]; // @[loaf.scala 276:58]
  assign _T_545 = _T_543[31:16]; // @[loaf.scala 276:58]
  assign _T_554 = AE_5_0__T_552_data;
  assign _T_555 = _T_554[15:0]; // @[loaf.scala 276:58]
  assign _T_556 = _T_554[31:16]; // @[loaf.scala 276:58]
  assign _T_565 = AE_6_0__T_563_data;
  assign _T_566 = _T_565[15:0]; // @[loaf.scala 276:58]
  assign _T_567 = _T_565[31:16]; // @[loaf.scala 276:58]
  assign _T_576 = AE_7_0__T_574_data;
  assign _T_577 = _T_576[15:0]; // @[loaf.scala 276:58]
  assign _T_578 = _T_576[31:16]; // @[loaf.scala 276:58]
  assign _T_587 = AE_0_1__T_585_data;
  assign _T_588 = _T_587[15:0]; // @[loaf.scala 276:58]
  assign _T_589 = _T_587[31:16]; // @[loaf.scala 276:58]
  assign _T_598 = AE_1_1__T_596_data;
  assign _T_599 = _T_598[15:0]; // @[loaf.scala 276:58]
  assign _T_600 = _T_598[31:16]; // @[loaf.scala 276:58]
  assign _T_609 = AE_2_1__T_607_data;
  assign _T_610 = _T_609[15:0]; // @[loaf.scala 276:58]
  assign _T_611 = _T_609[31:16]; // @[loaf.scala 276:58]
  assign _T_620 = AE_3_1__T_618_data;
  assign _T_621 = _T_620[15:0]; // @[loaf.scala 276:58]
  assign _T_622 = _T_620[31:16]; // @[loaf.scala 276:58]
  assign _T_631 = AE_4_1__T_629_data;
  assign _T_632 = _T_631[15:0]; // @[loaf.scala 276:58]
  assign _T_633 = _T_631[31:16]; // @[loaf.scala 276:58]
  assign _T_642 = AE_5_1__T_640_data;
  assign _T_643 = _T_642[15:0]; // @[loaf.scala 276:58]
  assign _T_644 = _T_642[31:16]; // @[loaf.scala 276:58]
  assign _T_653 = AE_6_1__T_651_data;
  assign _T_654 = _T_653[15:0]; // @[loaf.scala 276:58]
  assign _T_655 = _T_653[31:16]; // @[loaf.scala 276:58]
  assign _T_664 = AE_7_1__T_662_data;
  assign _T_665 = _T_664[15:0]; // @[loaf.scala 276:58]
  assign _T_666 = _T_664[31:16]; // @[loaf.scala 276:58]
  assign _T_675 = AE_0_2__T_673_data;
  assign _T_676 = _T_675[15:0]; // @[loaf.scala 276:58]
  assign _T_677 = _T_675[31:16]; // @[loaf.scala 276:58]
  assign _T_686 = AE_1_2__T_684_data;
  assign _T_687 = _T_686[15:0]; // @[loaf.scala 276:58]
  assign _T_688 = _T_686[31:16]; // @[loaf.scala 276:58]
  assign _T_697 = AE_2_2__T_695_data;
  assign _T_698 = _T_697[15:0]; // @[loaf.scala 276:58]
  assign _T_699 = _T_697[31:16]; // @[loaf.scala 276:58]
  assign _T_708 = AE_3_2__T_706_data;
  assign _T_709 = _T_708[15:0]; // @[loaf.scala 276:58]
  assign _T_710 = _T_708[31:16]; // @[loaf.scala 276:58]
  assign _T_719 = AE_4_2__T_717_data;
  assign _T_720 = _T_719[15:0]; // @[loaf.scala 276:58]
  assign _T_721 = _T_719[31:16]; // @[loaf.scala 276:58]
  assign _T_730 = AE_5_2__T_728_data;
  assign _T_731 = _T_730[15:0]; // @[loaf.scala 276:58]
  assign _T_732 = _T_730[31:16]; // @[loaf.scala 276:58]
  assign _T_741 = AE_6_2__T_739_data;
  assign _T_742 = _T_741[15:0]; // @[loaf.scala 276:58]
  assign _T_743 = _T_741[31:16]; // @[loaf.scala 276:58]
  assign _T_752 = AE_7_2__T_750_data;
  assign _T_753 = _T_752[15:0]; // @[loaf.scala 276:58]
  assign _T_754 = _T_752[31:16]; // @[loaf.scala 276:58]
  assign _T_763 = AE_0_3__T_761_data;
  assign _T_764 = _T_763[15:0]; // @[loaf.scala 276:58]
  assign _T_765 = _T_763[31:16]; // @[loaf.scala 276:58]
  assign _T_774 = AE_1_3__T_772_data;
  assign _T_775 = _T_774[15:0]; // @[loaf.scala 276:58]
  assign _T_776 = _T_774[31:16]; // @[loaf.scala 276:58]
  assign _T_785 = AE_2_3__T_783_data;
  assign _T_786 = _T_785[15:0]; // @[loaf.scala 276:58]
  assign _T_787 = _T_785[31:16]; // @[loaf.scala 276:58]
  assign _T_796 = AE_3_3__T_794_data;
  assign _T_797 = _T_796[15:0]; // @[loaf.scala 276:58]
  assign _T_798 = _T_796[31:16]; // @[loaf.scala 276:58]
  assign _T_807 = AE_4_3__T_805_data;
  assign _T_808 = _T_807[15:0]; // @[loaf.scala 276:58]
  assign _T_809 = _T_807[31:16]; // @[loaf.scala 276:58]
  assign _T_818 = AE_5_3__T_816_data;
  assign _T_819 = _T_818[15:0]; // @[loaf.scala 276:58]
  assign _T_820 = _T_818[31:16]; // @[loaf.scala 276:58]
  assign _T_829 = AE_6_3__T_827_data;
  assign _T_830 = _T_829[15:0]; // @[loaf.scala 276:58]
  assign _T_831 = _T_829[31:16]; // @[loaf.scala 276:58]
  assign _T_840 = AE_7_3__T_838_data;
  assign _T_841 = _T_840[15:0]; // @[loaf.scala 276:58]
  assign _T_842 = _T_840[31:16]; // @[loaf.scala 276:58]
  assign _T_851 = AE_0_4__T_849_data;
  assign _T_852 = _T_851[15:0]; // @[loaf.scala 276:58]
  assign _T_853 = _T_851[31:16]; // @[loaf.scala 276:58]
  assign _T_862 = AE_1_4__T_860_data;
  assign _T_863 = _T_862[15:0]; // @[loaf.scala 276:58]
  assign _T_864 = _T_862[31:16]; // @[loaf.scala 276:58]
  assign _T_873 = AE_2_4__T_871_data;
  assign _T_874 = _T_873[15:0]; // @[loaf.scala 276:58]
  assign _T_875 = _T_873[31:16]; // @[loaf.scala 276:58]
  assign _T_884 = AE_3_4__T_882_data;
  assign _T_885 = _T_884[15:0]; // @[loaf.scala 276:58]
  assign _T_886 = _T_884[31:16]; // @[loaf.scala 276:58]
  assign _T_895 = AE_4_4__T_893_data;
  assign _T_896 = _T_895[15:0]; // @[loaf.scala 276:58]
  assign _T_897 = _T_895[31:16]; // @[loaf.scala 276:58]
  assign _T_906 = AE_5_4__T_904_data;
  assign _T_907 = _T_906[15:0]; // @[loaf.scala 276:58]
  assign _T_908 = _T_906[31:16]; // @[loaf.scala 276:58]
  assign _T_917 = AE_6_4__T_915_data;
  assign _T_918 = _T_917[15:0]; // @[loaf.scala 276:58]
  assign _T_919 = _T_917[31:16]; // @[loaf.scala 276:58]
  assign _T_928 = AE_7_4__T_926_data;
  assign _T_929 = _T_928[15:0]; // @[loaf.scala 276:58]
  assign _T_930 = _T_928[31:16]; // @[loaf.scala 276:58]
  assign _T_939 = AE_0_5__T_937_data;
  assign _T_940 = _T_939[15:0]; // @[loaf.scala 276:58]
  assign _T_941 = _T_939[31:16]; // @[loaf.scala 276:58]
  assign _T_950 = AE_1_5__T_948_data;
  assign _T_951 = _T_950[15:0]; // @[loaf.scala 276:58]
  assign _T_952 = _T_950[31:16]; // @[loaf.scala 276:58]
  assign _T_961 = AE_2_5__T_959_data;
  assign _T_962 = _T_961[15:0]; // @[loaf.scala 276:58]
  assign _T_963 = _T_961[31:16]; // @[loaf.scala 276:58]
  assign _T_972 = AE_3_5__T_970_data;
  assign _T_973 = _T_972[15:0]; // @[loaf.scala 276:58]
  assign _T_974 = _T_972[31:16]; // @[loaf.scala 276:58]
  assign _T_983 = AE_4_5__T_981_data;
  assign _T_984 = _T_983[15:0]; // @[loaf.scala 276:58]
  assign _T_985 = _T_983[31:16]; // @[loaf.scala 276:58]
  assign _T_994 = AE_5_5__T_992_data;
  assign _T_995 = _T_994[15:0]; // @[loaf.scala 276:58]
  assign _T_996 = _T_994[31:16]; // @[loaf.scala 276:58]
  assign _T_1005 = AE_6_5__T_1003_data;
  assign _T_1006 = _T_1005[15:0]; // @[loaf.scala 276:58]
  assign _T_1007 = _T_1005[31:16]; // @[loaf.scala 276:58]
  assign _T_1016 = AE_7_5__T_1014_data;
  assign _T_1017 = _T_1016[15:0]; // @[loaf.scala 276:58]
  assign _T_1018 = _T_1016[31:16]; // @[loaf.scala 276:58]
  assign _T_1027 = AE_0_6__T_1025_data;
  assign _T_1028 = _T_1027[15:0]; // @[loaf.scala 276:58]
  assign _T_1029 = _T_1027[31:16]; // @[loaf.scala 276:58]
  assign _T_1038 = AE_1_6__T_1036_data;
  assign _T_1039 = _T_1038[15:0]; // @[loaf.scala 276:58]
  assign _T_1040 = _T_1038[31:16]; // @[loaf.scala 276:58]
  assign _T_1049 = AE_2_6__T_1047_data;
  assign _T_1050 = _T_1049[15:0]; // @[loaf.scala 276:58]
  assign _T_1051 = _T_1049[31:16]; // @[loaf.scala 276:58]
  assign _T_1060 = AE_3_6__T_1058_data;
  assign _T_1061 = _T_1060[15:0]; // @[loaf.scala 276:58]
  assign _T_1062 = _T_1060[31:16]; // @[loaf.scala 276:58]
  assign _T_1071 = AE_4_6__T_1069_data;
  assign _T_1072 = _T_1071[15:0]; // @[loaf.scala 276:58]
  assign _T_1073 = _T_1071[31:16]; // @[loaf.scala 276:58]
  assign _T_1082 = AE_5_6__T_1080_data;
  assign _T_1083 = _T_1082[15:0]; // @[loaf.scala 276:58]
  assign _T_1084 = _T_1082[31:16]; // @[loaf.scala 276:58]
  assign _T_1093 = AE_6_6__T_1091_data;
  assign _T_1094 = _T_1093[15:0]; // @[loaf.scala 276:58]
  assign _T_1095 = _T_1093[31:16]; // @[loaf.scala 276:58]
  assign _T_1104 = AE_7_6__T_1102_data;
  assign _T_1105 = _T_1104[15:0]; // @[loaf.scala 276:58]
  assign _T_1106 = _T_1104[31:16]; // @[loaf.scala 276:58]
  assign _T_1115 = AE_0_7__T_1113_data;
  assign _T_1116 = _T_1115[15:0]; // @[loaf.scala 276:58]
  assign _T_1117 = _T_1115[31:16]; // @[loaf.scala 276:58]
  assign _T_1126 = AE_1_7__T_1124_data;
  assign _T_1127 = _T_1126[15:0]; // @[loaf.scala 276:58]
  assign _T_1128 = _T_1126[31:16]; // @[loaf.scala 276:58]
  assign _T_1137 = AE_2_7__T_1135_data;
  assign _T_1138 = _T_1137[15:0]; // @[loaf.scala 276:58]
  assign _T_1139 = _T_1137[31:16]; // @[loaf.scala 276:58]
  assign _T_1148 = AE_3_7__T_1146_data;
  assign _T_1149 = _T_1148[15:0]; // @[loaf.scala 276:58]
  assign _T_1150 = _T_1148[31:16]; // @[loaf.scala 276:58]
  assign _T_1159 = AE_4_7__T_1157_data;
  assign _T_1160 = _T_1159[15:0]; // @[loaf.scala 276:58]
  assign _T_1161 = _T_1159[31:16]; // @[loaf.scala 276:58]
  assign _T_1170 = AE_5_7__T_1168_data;
  assign _T_1171 = _T_1170[15:0]; // @[loaf.scala 276:58]
  assign _T_1172 = _T_1170[31:16]; // @[loaf.scala 276:58]
  assign _T_1181 = AE_6_7__T_1179_data;
  assign _T_1182 = _T_1181[15:0]; // @[loaf.scala 276:58]
  assign _T_1183 = _T_1181[31:16]; // @[loaf.scala 276:58]
  assign _T_1192 = AE_7_7__T_1190_data;
  assign _T_1193 = _T_1192[15:0]; // @[loaf.scala 276:58]
  assign _T_1194 = _T_1192[31:16]; // @[loaf.scala 276:58]
  assign _T_1196 = BFbuf_e > AEbuf_0_0_e; // @[loaf.scala 292:22]
  assign _T_1198 = AEbuf_0_0_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_1200 = AEbuf_0_0_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_1202 = BFbuf_a - AEbuf_0_0_a; // @[loaf.scala 295:34]
  assign _T_1204 = ab2_0_0 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2003 = _T_1204 ? 16'hcc : ab2_0_0; // @[loaf.scala 298:37]
  assign _T_1205 = {$signed(o2_0), 10'h0}; // @[loaf.scala 302:38]
  assign _T_1206 = macs_0_0_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_1208 = BFbuf_e > AEbuf_1_0_e; // @[loaf.scala 292:22]
  assign _T_1210 = AEbuf_1_0_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_1212 = AEbuf_1_0_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_1214 = BFbuf_a - AEbuf_1_0_a; // @[loaf.scala 295:34]
  assign _T_1216 = ab2_1_0 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2006 = _T_1216 ? 16'hcc : ab2_1_0; // @[loaf.scala 298:37]
  assign _T_1217 = {$signed(o2_1), 10'h0}; // @[loaf.scala 302:38]
  assign _T_1218 = macs_1_0_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_1220 = BFbuf_e > AEbuf_2_0_e; // @[loaf.scala 292:22]
  assign _T_1222 = AEbuf_2_0_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_1224 = AEbuf_2_0_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_1226 = BFbuf_a - AEbuf_2_0_a; // @[loaf.scala 295:34]
  assign _T_1228 = ab2_2_0 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2009 = _T_1228 ? 16'hcc : ab2_2_0; // @[loaf.scala 298:37]
  assign _T_1229 = {$signed(o2_2), 10'h0}; // @[loaf.scala 302:38]
  assign _T_1230 = macs_2_0_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_1232 = BFbuf_e > AEbuf_3_0_e; // @[loaf.scala 292:22]
  assign _T_1234 = AEbuf_3_0_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_1236 = AEbuf_3_0_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_1238 = BFbuf_a - AEbuf_3_0_a; // @[loaf.scala 295:34]
  assign _T_1240 = ab2_3_0 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2012 = _T_1240 ? 16'hcc : ab2_3_0; // @[loaf.scala 298:37]
  assign _T_1241 = {$signed(o2_3), 10'h0}; // @[loaf.scala 302:38]
  assign _T_1242 = macs_3_0_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_1244 = BFbuf_e > AEbuf_4_0_e; // @[loaf.scala 292:22]
  assign _T_1246 = AEbuf_4_0_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_1248 = AEbuf_4_0_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_1250 = BFbuf_a - AEbuf_4_0_a; // @[loaf.scala 295:34]
  assign _T_1252 = ab2_4_0 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2015 = _T_1252 ? 16'hcc : ab2_4_0; // @[loaf.scala 298:37]
  assign _T_1253 = {$signed(o2_4), 10'h0}; // @[loaf.scala 302:38]
  assign _T_1254 = macs_4_0_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_1256 = BFbuf_e > AEbuf_5_0_e; // @[loaf.scala 292:22]
  assign _T_1258 = AEbuf_5_0_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_1260 = AEbuf_5_0_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_1262 = BFbuf_a - AEbuf_5_0_a; // @[loaf.scala 295:34]
  assign _T_1264 = ab2_5_0 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2018 = _T_1264 ? 16'hcc : ab2_5_0; // @[loaf.scala 298:37]
  assign _T_1265 = {$signed(o2_5), 10'h0}; // @[loaf.scala 302:38]
  assign _T_1266 = macs_5_0_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_1268 = BFbuf_e > AEbuf_6_0_e; // @[loaf.scala 292:22]
  assign _T_1270 = AEbuf_6_0_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_1272 = AEbuf_6_0_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_1274 = BFbuf_a - AEbuf_6_0_a; // @[loaf.scala 295:34]
  assign _T_1276 = ab2_6_0 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2021 = _T_1276 ? 16'hcc : ab2_6_0; // @[loaf.scala 298:37]
  assign _T_1277 = {$signed(o2_6), 10'h0}; // @[loaf.scala 302:38]
  assign _T_1278 = macs_6_0_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_1280 = BFbuf_e > AEbuf_7_0_e; // @[loaf.scala 292:22]
  assign _T_1282 = AEbuf_7_0_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_1284 = AEbuf_7_0_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_1286 = BFbuf_a - AEbuf_7_0_a; // @[loaf.scala 295:34]
  assign _T_1288 = ab2_7_0 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2024 = _T_1288 ? 16'hcc : ab2_7_0; // @[loaf.scala 298:37]
  assign _T_1289 = {$signed(o2_7), 10'h0}; // @[loaf.scala 302:38]
  assign _T_1290 = macs_7_0_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_1292 = $signed(_T_1206) < $signed(_T_1218); // @[loaf.scala 327:24]
  assign _GEN_2025 = _T_1292 ? $signed(_T_1206) : $signed(_T_1218); // @[loaf.scala 327:29]
  assign _T_1294 = $signed(_T_1230) < $signed(_T_1242); // @[loaf.scala 327:24]
  assign _GEN_2026 = _T_1294 ? $signed(_T_1230) : $signed(_T_1242); // @[loaf.scala 327:29]
  assign _T_1296 = $signed(_T_1254) < $signed(_T_1266); // @[loaf.scala 327:24]
  assign _GEN_2027 = _T_1296 ? $signed(_T_1254) : $signed(_T_1266); // @[loaf.scala 327:29]
  assign _T_1298 = $signed(_T_1278) < $signed(_T_1290); // @[loaf.scala 327:24]
  assign _GEN_2028 = _T_1298 ? $signed(_T_1278) : $signed(_T_1290); // @[loaf.scala 327:29]
  assign _T_1300 = $signed(tm8_0_0) < $signed(tm8_1_0); // @[loaf.scala 327:24]
  assign _T_1302 = $signed(tm8_2_0) < $signed(tm8_3_0); // @[loaf.scala 327:24]
  assign _T_1304 = $signed(tm9_0_0) < $signed(tm9_1_0); // @[loaf.scala 327:24]
  assign _T_1306 = $signed(tmc_0_0) < $signed(best_0); // @[loaf.scala 354:43]
  assign _T_1307 = _T_448 | _T_1306; // @[loaf.scala 354:35]
  assign _T_1309 = BFbuf_e > AEbuf_0_1_e; // @[loaf.scala 292:22]
  assign _T_1311 = AEbuf_0_1_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_1313 = AEbuf_0_1_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_1315 = BFbuf_a - AEbuf_0_1_a; // @[loaf.scala 295:34]
  assign _T_1317 = ab2_0_1 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2035 = _T_1317 ? 16'hcc : ab2_0_1; // @[loaf.scala 298:37]
  assign _T_1319 = macs_0_1_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_1321 = BFbuf_e > AEbuf_1_1_e; // @[loaf.scala 292:22]
  assign _T_1323 = AEbuf_1_1_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_1325 = AEbuf_1_1_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_1327 = BFbuf_a - AEbuf_1_1_a; // @[loaf.scala 295:34]
  assign _T_1329 = ab2_1_1 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2038 = _T_1329 ? 16'hcc : ab2_1_1; // @[loaf.scala 298:37]
  assign _T_1331 = macs_1_1_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_1333 = BFbuf_e > AEbuf_2_1_e; // @[loaf.scala 292:22]
  assign _T_1335 = AEbuf_2_1_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_1337 = AEbuf_2_1_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_1339 = BFbuf_a - AEbuf_2_1_a; // @[loaf.scala 295:34]
  assign _T_1341 = ab2_2_1 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2041 = _T_1341 ? 16'hcc : ab2_2_1; // @[loaf.scala 298:37]
  assign _T_1343 = macs_2_1_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_1345 = BFbuf_e > AEbuf_3_1_e; // @[loaf.scala 292:22]
  assign _T_1347 = AEbuf_3_1_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_1349 = AEbuf_3_1_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_1351 = BFbuf_a - AEbuf_3_1_a; // @[loaf.scala 295:34]
  assign _T_1353 = ab2_3_1 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2044 = _T_1353 ? 16'hcc : ab2_3_1; // @[loaf.scala 298:37]
  assign _T_1355 = macs_3_1_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_1357 = BFbuf_e > AEbuf_4_1_e; // @[loaf.scala 292:22]
  assign _T_1359 = AEbuf_4_1_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_1361 = AEbuf_4_1_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_1363 = BFbuf_a - AEbuf_4_1_a; // @[loaf.scala 295:34]
  assign _T_1365 = ab2_4_1 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2047 = _T_1365 ? 16'hcc : ab2_4_1; // @[loaf.scala 298:37]
  assign _T_1367 = macs_4_1_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_1369 = BFbuf_e > AEbuf_5_1_e; // @[loaf.scala 292:22]
  assign _T_1371 = AEbuf_5_1_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_1373 = AEbuf_5_1_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_1375 = BFbuf_a - AEbuf_5_1_a; // @[loaf.scala 295:34]
  assign _T_1377 = ab2_5_1 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2050 = _T_1377 ? 16'hcc : ab2_5_1; // @[loaf.scala 298:37]
  assign _T_1379 = macs_5_1_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_1381 = BFbuf_e > AEbuf_6_1_e; // @[loaf.scala 292:22]
  assign _T_1383 = AEbuf_6_1_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_1385 = AEbuf_6_1_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_1387 = BFbuf_a - AEbuf_6_1_a; // @[loaf.scala 295:34]
  assign _T_1389 = ab2_6_1 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2053 = _T_1389 ? 16'hcc : ab2_6_1; // @[loaf.scala 298:37]
  assign _T_1391 = macs_6_1_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_1393 = BFbuf_e > AEbuf_7_1_e; // @[loaf.scala 292:22]
  assign _T_1395 = AEbuf_7_1_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_1397 = AEbuf_7_1_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_1399 = BFbuf_a - AEbuf_7_1_a; // @[loaf.scala 295:34]
  assign _T_1401 = ab2_7_1 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2056 = _T_1401 ? 16'hcc : ab2_7_1; // @[loaf.scala 298:37]
  assign _T_1403 = macs_7_1_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_1405 = $signed(_T_1319) < $signed(_T_1331); // @[loaf.scala 327:24]
  assign _GEN_2057 = _T_1405 ? $signed(_T_1319) : $signed(_T_1331); // @[loaf.scala 327:29]
  assign _T_1407 = $signed(_T_1343) < $signed(_T_1355); // @[loaf.scala 327:24]
  assign _GEN_2058 = _T_1407 ? $signed(_T_1343) : $signed(_T_1355); // @[loaf.scala 327:29]
  assign _T_1409 = $signed(_T_1367) < $signed(_T_1379); // @[loaf.scala 327:24]
  assign _GEN_2059 = _T_1409 ? $signed(_T_1367) : $signed(_T_1379); // @[loaf.scala 327:29]
  assign _T_1411 = $signed(_T_1391) < $signed(_T_1403); // @[loaf.scala 327:24]
  assign _GEN_2060 = _T_1411 ? $signed(_T_1391) : $signed(_T_1403); // @[loaf.scala 327:29]
  assign _T_1413 = $signed(tm8_0_1) < $signed(tm8_1_1); // @[loaf.scala 327:24]
  assign _T_1415 = $signed(tm8_2_1) < $signed(tm8_3_1); // @[loaf.scala 327:24]
  assign _T_1417 = $signed(tm9_0_1) < $signed(tm9_1_1); // @[loaf.scala 327:24]
  assign _T_1419 = $signed(tmc_0_1) < $signed(best_1); // @[loaf.scala 354:43]
  assign _T_1420 = _T_448 | _T_1419; // @[loaf.scala 354:35]
  assign _T_1422 = BFbuf_e > AEbuf_0_2_e; // @[loaf.scala 292:22]
  assign _T_1424 = AEbuf_0_2_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_1426 = AEbuf_0_2_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_1428 = BFbuf_a - AEbuf_0_2_a; // @[loaf.scala 295:34]
  assign _T_1430 = ab2_0_2 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2067 = _T_1430 ? 16'hcc : ab2_0_2; // @[loaf.scala 298:37]
  assign _T_1432 = macs_0_2_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_1434 = BFbuf_e > AEbuf_1_2_e; // @[loaf.scala 292:22]
  assign _T_1436 = AEbuf_1_2_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_1438 = AEbuf_1_2_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_1440 = BFbuf_a - AEbuf_1_2_a; // @[loaf.scala 295:34]
  assign _T_1442 = ab2_1_2 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2070 = _T_1442 ? 16'hcc : ab2_1_2; // @[loaf.scala 298:37]
  assign _T_1444 = macs_1_2_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_1446 = BFbuf_e > AEbuf_2_2_e; // @[loaf.scala 292:22]
  assign _T_1448 = AEbuf_2_2_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_1450 = AEbuf_2_2_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_1452 = BFbuf_a - AEbuf_2_2_a; // @[loaf.scala 295:34]
  assign _T_1454 = ab2_2_2 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2073 = _T_1454 ? 16'hcc : ab2_2_2; // @[loaf.scala 298:37]
  assign _T_1456 = macs_2_2_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_1458 = BFbuf_e > AEbuf_3_2_e; // @[loaf.scala 292:22]
  assign _T_1460 = AEbuf_3_2_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_1462 = AEbuf_3_2_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_1464 = BFbuf_a - AEbuf_3_2_a; // @[loaf.scala 295:34]
  assign _T_1466 = ab2_3_2 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2076 = _T_1466 ? 16'hcc : ab2_3_2; // @[loaf.scala 298:37]
  assign _T_1468 = macs_3_2_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_1470 = BFbuf_e > AEbuf_4_2_e; // @[loaf.scala 292:22]
  assign _T_1472 = AEbuf_4_2_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_1474 = AEbuf_4_2_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_1476 = BFbuf_a - AEbuf_4_2_a; // @[loaf.scala 295:34]
  assign _T_1478 = ab2_4_2 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2079 = _T_1478 ? 16'hcc : ab2_4_2; // @[loaf.scala 298:37]
  assign _T_1480 = macs_4_2_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_1482 = BFbuf_e > AEbuf_5_2_e; // @[loaf.scala 292:22]
  assign _T_1484 = AEbuf_5_2_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_1486 = AEbuf_5_2_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_1488 = BFbuf_a - AEbuf_5_2_a; // @[loaf.scala 295:34]
  assign _T_1490 = ab2_5_2 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2082 = _T_1490 ? 16'hcc : ab2_5_2; // @[loaf.scala 298:37]
  assign _T_1492 = macs_5_2_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_1494 = BFbuf_e > AEbuf_6_2_e; // @[loaf.scala 292:22]
  assign _T_1496 = AEbuf_6_2_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_1498 = AEbuf_6_2_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_1500 = BFbuf_a - AEbuf_6_2_a; // @[loaf.scala 295:34]
  assign _T_1502 = ab2_6_2 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2085 = _T_1502 ? 16'hcc : ab2_6_2; // @[loaf.scala 298:37]
  assign _T_1504 = macs_6_2_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_1506 = BFbuf_e > AEbuf_7_2_e; // @[loaf.scala 292:22]
  assign _T_1508 = AEbuf_7_2_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_1510 = AEbuf_7_2_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_1512 = BFbuf_a - AEbuf_7_2_a; // @[loaf.scala 295:34]
  assign _T_1514 = ab2_7_2 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2088 = _T_1514 ? 16'hcc : ab2_7_2; // @[loaf.scala 298:37]
  assign _T_1516 = macs_7_2_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_1518 = $signed(_T_1432) < $signed(_T_1444); // @[loaf.scala 327:24]
  assign _GEN_2089 = _T_1518 ? $signed(_T_1432) : $signed(_T_1444); // @[loaf.scala 327:29]
  assign _T_1520 = $signed(_T_1456) < $signed(_T_1468); // @[loaf.scala 327:24]
  assign _GEN_2090 = _T_1520 ? $signed(_T_1456) : $signed(_T_1468); // @[loaf.scala 327:29]
  assign _T_1522 = $signed(_T_1480) < $signed(_T_1492); // @[loaf.scala 327:24]
  assign _GEN_2091 = _T_1522 ? $signed(_T_1480) : $signed(_T_1492); // @[loaf.scala 327:29]
  assign _T_1524 = $signed(_T_1504) < $signed(_T_1516); // @[loaf.scala 327:24]
  assign _GEN_2092 = _T_1524 ? $signed(_T_1504) : $signed(_T_1516); // @[loaf.scala 327:29]
  assign _T_1526 = $signed(tm8_0_2) < $signed(tm8_1_2); // @[loaf.scala 327:24]
  assign _T_1528 = $signed(tm8_2_2) < $signed(tm8_3_2); // @[loaf.scala 327:24]
  assign _T_1530 = $signed(tm9_0_2) < $signed(tm9_1_2); // @[loaf.scala 327:24]
  assign _T_1532 = $signed(tmc_0_2) < $signed(best_2); // @[loaf.scala 354:43]
  assign _T_1533 = _T_448 | _T_1532; // @[loaf.scala 354:35]
  assign _T_1535 = BFbuf_e > AEbuf_0_3_e; // @[loaf.scala 292:22]
  assign _T_1537 = AEbuf_0_3_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_1539 = AEbuf_0_3_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_1541 = BFbuf_a - AEbuf_0_3_a; // @[loaf.scala 295:34]
  assign _T_1543 = ab2_0_3 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2099 = _T_1543 ? 16'hcc : ab2_0_3; // @[loaf.scala 298:37]
  assign _T_1545 = macs_0_3_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_1547 = BFbuf_e > AEbuf_1_3_e; // @[loaf.scala 292:22]
  assign _T_1549 = AEbuf_1_3_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_1551 = AEbuf_1_3_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_1553 = BFbuf_a - AEbuf_1_3_a; // @[loaf.scala 295:34]
  assign _T_1555 = ab2_1_3 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2102 = _T_1555 ? 16'hcc : ab2_1_3; // @[loaf.scala 298:37]
  assign _T_1557 = macs_1_3_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_1559 = BFbuf_e > AEbuf_2_3_e; // @[loaf.scala 292:22]
  assign _T_1561 = AEbuf_2_3_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_1563 = AEbuf_2_3_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_1565 = BFbuf_a - AEbuf_2_3_a; // @[loaf.scala 295:34]
  assign _T_1567 = ab2_2_3 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2105 = _T_1567 ? 16'hcc : ab2_2_3; // @[loaf.scala 298:37]
  assign _T_1569 = macs_2_3_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_1571 = BFbuf_e > AEbuf_3_3_e; // @[loaf.scala 292:22]
  assign _T_1573 = AEbuf_3_3_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_1575 = AEbuf_3_3_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_1577 = BFbuf_a - AEbuf_3_3_a; // @[loaf.scala 295:34]
  assign _T_1579 = ab2_3_3 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2108 = _T_1579 ? 16'hcc : ab2_3_3; // @[loaf.scala 298:37]
  assign _T_1581 = macs_3_3_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_1583 = BFbuf_e > AEbuf_4_3_e; // @[loaf.scala 292:22]
  assign _T_1585 = AEbuf_4_3_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_1587 = AEbuf_4_3_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_1589 = BFbuf_a - AEbuf_4_3_a; // @[loaf.scala 295:34]
  assign _T_1591 = ab2_4_3 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2111 = _T_1591 ? 16'hcc : ab2_4_3; // @[loaf.scala 298:37]
  assign _T_1593 = macs_4_3_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_1595 = BFbuf_e > AEbuf_5_3_e; // @[loaf.scala 292:22]
  assign _T_1597 = AEbuf_5_3_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_1599 = AEbuf_5_3_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_1601 = BFbuf_a - AEbuf_5_3_a; // @[loaf.scala 295:34]
  assign _T_1603 = ab2_5_3 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2114 = _T_1603 ? 16'hcc : ab2_5_3; // @[loaf.scala 298:37]
  assign _T_1605 = macs_5_3_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_1607 = BFbuf_e > AEbuf_6_3_e; // @[loaf.scala 292:22]
  assign _T_1609 = AEbuf_6_3_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_1611 = AEbuf_6_3_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_1613 = BFbuf_a - AEbuf_6_3_a; // @[loaf.scala 295:34]
  assign _T_1615 = ab2_6_3 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2117 = _T_1615 ? 16'hcc : ab2_6_3; // @[loaf.scala 298:37]
  assign _T_1617 = macs_6_3_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_1619 = BFbuf_e > AEbuf_7_3_e; // @[loaf.scala 292:22]
  assign _T_1621 = AEbuf_7_3_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_1623 = AEbuf_7_3_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_1625 = BFbuf_a - AEbuf_7_3_a; // @[loaf.scala 295:34]
  assign _T_1627 = ab2_7_3 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2120 = _T_1627 ? 16'hcc : ab2_7_3; // @[loaf.scala 298:37]
  assign _T_1629 = macs_7_3_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_1631 = $signed(_T_1545) < $signed(_T_1557); // @[loaf.scala 327:24]
  assign _GEN_2121 = _T_1631 ? $signed(_T_1545) : $signed(_T_1557); // @[loaf.scala 327:29]
  assign _T_1633 = $signed(_T_1569) < $signed(_T_1581); // @[loaf.scala 327:24]
  assign _GEN_2122 = _T_1633 ? $signed(_T_1569) : $signed(_T_1581); // @[loaf.scala 327:29]
  assign _T_1635 = $signed(_T_1593) < $signed(_T_1605); // @[loaf.scala 327:24]
  assign _GEN_2123 = _T_1635 ? $signed(_T_1593) : $signed(_T_1605); // @[loaf.scala 327:29]
  assign _T_1637 = $signed(_T_1617) < $signed(_T_1629); // @[loaf.scala 327:24]
  assign _GEN_2124 = _T_1637 ? $signed(_T_1617) : $signed(_T_1629); // @[loaf.scala 327:29]
  assign _T_1639 = $signed(tm8_0_3) < $signed(tm8_1_3); // @[loaf.scala 327:24]
  assign _T_1641 = $signed(tm8_2_3) < $signed(tm8_3_3); // @[loaf.scala 327:24]
  assign _T_1643 = $signed(tm9_0_3) < $signed(tm9_1_3); // @[loaf.scala 327:24]
  assign _T_1645 = $signed(tmc_0_3) < $signed(best_3); // @[loaf.scala 354:43]
  assign _T_1646 = _T_448 | _T_1645; // @[loaf.scala 354:35]
  assign _T_1648 = BFbuf_e > AEbuf_0_4_e; // @[loaf.scala 292:22]
  assign _T_1650 = AEbuf_0_4_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_1652 = AEbuf_0_4_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_1654 = BFbuf_a - AEbuf_0_4_a; // @[loaf.scala 295:34]
  assign _T_1656 = ab2_0_4 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2131 = _T_1656 ? 16'hcc : ab2_0_4; // @[loaf.scala 298:37]
  assign _T_1658 = macs_0_4_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_1660 = BFbuf_e > AEbuf_1_4_e; // @[loaf.scala 292:22]
  assign _T_1662 = AEbuf_1_4_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_1664 = AEbuf_1_4_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_1666 = BFbuf_a - AEbuf_1_4_a; // @[loaf.scala 295:34]
  assign _T_1668 = ab2_1_4 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2134 = _T_1668 ? 16'hcc : ab2_1_4; // @[loaf.scala 298:37]
  assign _T_1670 = macs_1_4_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_1672 = BFbuf_e > AEbuf_2_4_e; // @[loaf.scala 292:22]
  assign _T_1674 = AEbuf_2_4_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_1676 = AEbuf_2_4_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_1678 = BFbuf_a - AEbuf_2_4_a; // @[loaf.scala 295:34]
  assign _T_1680 = ab2_2_4 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2137 = _T_1680 ? 16'hcc : ab2_2_4; // @[loaf.scala 298:37]
  assign _T_1682 = macs_2_4_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_1684 = BFbuf_e > AEbuf_3_4_e; // @[loaf.scala 292:22]
  assign _T_1686 = AEbuf_3_4_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_1688 = AEbuf_3_4_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_1690 = BFbuf_a - AEbuf_3_4_a; // @[loaf.scala 295:34]
  assign _T_1692 = ab2_3_4 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2140 = _T_1692 ? 16'hcc : ab2_3_4; // @[loaf.scala 298:37]
  assign _T_1694 = macs_3_4_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_1696 = BFbuf_e > AEbuf_4_4_e; // @[loaf.scala 292:22]
  assign _T_1698 = AEbuf_4_4_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_1700 = AEbuf_4_4_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_1702 = BFbuf_a - AEbuf_4_4_a; // @[loaf.scala 295:34]
  assign _T_1704 = ab2_4_4 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2143 = _T_1704 ? 16'hcc : ab2_4_4; // @[loaf.scala 298:37]
  assign _T_1706 = macs_4_4_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_1708 = BFbuf_e > AEbuf_5_4_e; // @[loaf.scala 292:22]
  assign _T_1710 = AEbuf_5_4_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_1712 = AEbuf_5_4_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_1714 = BFbuf_a - AEbuf_5_4_a; // @[loaf.scala 295:34]
  assign _T_1716 = ab2_5_4 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2146 = _T_1716 ? 16'hcc : ab2_5_4; // @[loaf.scala 298:37]
  assign _T_1718 = macs_5_4_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_1720 = BFbuf_e > AEbuf_6_4_e; // @[loaf.scala 292:22]
  assign _T_1722 = AEbuf_6_4_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_1724 = AEbuf_6_4_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_1726 = BFbuf_a - AEbuf_6_4_a; // @[loaf.scala 295:34]
  assign _T_1728 = ab2_6_4 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2149 = _T_1728 ? 16'hcc : ab2_6_4; // @[loaf.scala 298:37]
  assign _T_1730 = macs_6_4_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_1732 = BFbuf_e > AEbuf_7_4_e; // @[loaf.scala 292:22]
  assign _T_1734 = AEbuf_7_4_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_1736 = AEbuf_7_4_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_1738 = BFbuf_a - AEbuf_7_4_a; // @[loaf.scala 295:34]
  assign _T_1740 = ab2_7_4 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2152 = _T_1740 ? 16'hcc : ab2_7_4; // @[loaf.scala 298:37]
  assign _T_1742 = macs_7_4_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_1744 = $signed(_T_1658) < $signed(_T_1670); // @[loaf.scala 327:24]
  assign _GEN_2153 = _T_1744 ? $signed(_T_1658) : $signed(_T_1670); // @[loaf.scala 327:29]
  assign _T_1746 = $signed(_T_1682) < $signed(_T_1694); // @[loaf.scala 327:24]
  assign _GEN_2154 = _T_1746 ? $signed(_T_1682) : $signed(_T_1694); // @[loaf.scala 327:29]
  assign _T_1748 = $signed(_T_1706) < $signed(_T_1718); // @[loaf.scala 327:24]
  assign _GEN_2155 = _T_1748 ? $signed(_T_1706) : $signed(_T_1718); // @[loaf.scala 327:29]
  assign _T_1750 = $signed(_T_1730) < $signed(_T_1742); // @[loaf.scala 327:24]
  assign _GEN_2156 = _T_1750 ? $signed(_T_1730) : $signed(_T_1742); // @[loaf.scala 327:29]
  assign _T_1752 = $signed(tm8_0_4) < $signed(tm8_1_4); // @[loaf.scala 327:24]
  assign _T_1754 = $signed(tm8_2_4) < $signed(tm8_3_4); // @[loaf.scala 327:24]
  assign _T_1756 = $signed(tm9_0_4) < $signed(tm9_1_4); // @[loaf.scala 327:24]
  assign _T_1758 = $signed(tmc_0_4) < $signed(best_4); // @[loaf.scala 354:43]
  assign _T_1759 = _T_448 | _T_1758; // @[loaf.scala 354:35]
  assign _T_1761 = BFbuf_e > AEbuf_0_5_e; // @[loaf.scala 292:22]
  assign _T_1763 = AEbuf_0_5_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_1765 = AEbuf_0_5_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_1767 = BFbuf_a - AEbuf_0_5_a; // @[loaf.scala 295:34]
  assign _T_1769 = ab2_0_5 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2163 = _T_1769 ? 16'hcc : ab2_0_5; // @[loaf.scala 298:37]
  assign _T_1771 = macs_0_5_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_1773 = BFbuf_e > AEbuf_1_5_e; // @[loaf.scala 292:22]
  assign _T_1775 = AEbuf_1_5_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_1777 = AEbuf_1_5_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_1779 = BFbuf_a - AEbuf_1_5_a; // @[loaf.scala 295:34]
  assign _T_1781 = ab2_1_5 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2166 = _T_1781 ? 16'hcc : ab2_1_5; // @[loaf.scala 298:37]
  assign _T_1783 = macs_1_5_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_1785 = BFbuf_e > AEbuf_2_5_e; // @[loaf.scala 292:22]
  assign _T_1787 = AEbuf_2_5_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_1789 = AEbuf_2_5_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_1791 = BFbuf_a - AEbuf_2_5_a; // @[loaf.scala 295:34]
  assign _T_1793 = ab2_2_5 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2169 = _T_1793 ? 16'hcc : ab2_2_5; // @[loaf.scala 298:37]
  assign _T_1795 = macs_2_5_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_1797 = BFbuf_e > AEbuf_3_5_e; // @[loaf.scala 292:22]
  assign _T_1799 = AEbuf_3_5_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_1801 = AEbuf_3_5_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_1803 = BFbuf_a - AEbuf_3_5_a; // @[loaf.scala 295:34]
  assign _T_1805 = ab2_3_5 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2172 = _T_1805 ? 16'hcc : ab2_3_5; // @[loaf.scala 298:37]
  assign _T_1807 = macs_3_5_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_1809 = BFbuf_e > AEbuf_4_5_e; // @[loaf.scala 292:22]
  assign _T_1811 = AEbuf_4_5_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_1813 = AEbuf_4_5_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_1815 = BFbuf_a - AEbuf_4_5_a; // @[loaf.scala 295:34]
  assign _T_1817 = ab2_4_5 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2175 = _T_1817 ? 16'hcc : ab2_4_5; // @[loaf.scala 298:37]
  assign _T_1819 = macs_4_5_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_1821 = BFbuf_e > AEbuf_5_5_e; // @[loaf.scala 292:22]
  assign _T_1823 = AEbuf_5_5_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_1825 = AEbuf_5_5_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_1827 = BFbuf_a - AEbuf_5_5_a; // @[loaf.scala 295:34]
  assign _T_1829 = ab2_5_5 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2178 = _T_1829 ? 16'hcc : ab2_5_5; // @[loaf.scala 298:37]
  assign _T_1831 = macs_5_5_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_1833 = BFbuf_e > AEbuf_6_5_e; // @[loaf.scala 292:22]
  assign _T_1835 = AEbuf_6_5_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_1837 = AEbuf_6_5_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_1839 = BFbuf_a - AEbuf_6_5_a; // @[loaf.scala 295:34]
  assign _T_1841 = ab2_6_5 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2181 = _T_1841 ? 16'hcc : ab2_6_5; // @[loaf.scala 298:37]
  assign _T_1843 = macs_6_5_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_1845 = BFbuf_e > AEbuf_7_5_e; // @[loaf.scala 292:22]
  assign _T_1847 = AEbuf_7_5_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_1849 = AEbuf_7_5_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_1851 = BFbuf_a - AEbuf_7_5_a; // @[loaf.scala 295:34]
  assign _T_1853 = ab2_7_5 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2184 = _T_1853 ? 16'hcc : ab2_7_5; // @[loaf.scala 298:37]
  assign _T_1855 = macs_7_5_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_1857 = $signed(_T_1771) < $signed(_T_1783); // @[loaf.scala 327:24]
  assign _GEN_2185 = _T_1857 ? $signed(_T_1771) : $signed(_T_1783); // @[loaf.scala 327:29]
  assign _T_1859 = $signed(_T_1795) < $signed(_T_1807); // @[loaf.scala 327:24]
  assign _GEN_2186 = _T_1859 ? $signed(_T_1795) : $signed(_T_1807); // @[loaf.scala 327:29]
  assign _T_1861 = $signed(_T_1819) < $signed(_T_1831); // @[loaf.scala 327:24]
  assign _GEN_2187 = _T_1861 ? $signed(_T_1819) : $signed(_T_1831); // @[loaf.scala 327:29]
  assign _T_1863 = $signed(_T_1843) < $signed(_T_1855); // @[loaf.scala 327:24]
  assign _GEN_2188 = _T_1863 ? $signed(_T_1843) : $signed(_T_1855); // @[loaf.scala 327:29]
  assign _T_1865 = $signed(tm8_0_5) < $signed(tm8_1_5); // @[loaf.scala 327:24]
  assign _T_1867 = $signed(tm8_2_5) < $signed(tm8_3_5); // @[loaf.scala 327:24]
  assign _T_1869 = $signed(tm9_0_5) < $signed(tm9_1_5); // @[loaf.scala 327:24]
  assign _T_1871 = $signed(tmc_0_5) < $signed(best_5); // @[loaf.scala 354:43]
  assign _T_1872 = _T_448 | _T_1871; // @[loaf.scala 354:35]
  assign _T_1874 = BFbuf_e > AEbuf_0_6_e; // @[loaf.scala 292:22]
  assign _T_1876 = AEbuf_0_6_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_1878 = AEbuf_0_6_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_1880 = BFbuf_a - AEbuf_0_6_a; // @[loaf.scala 295:34]
  assign _T_1882 = ab2_0_6 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2195 = _T_1882 ? 16'hcc : ab2_0_6; // @[loaf.scala 298:37]
  assign _T_1884 = macs_0_6_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_1886 = BFbuf_e > AEbuf_1_6_e; // @[loaf.scala 292:22]
  assign _T_1888 = AEbuf_1_6_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_1890 = AEbuf_1_6_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_1892 = BFbuf_a - AEbuf_1_6_a; // @[loaf.scala 295:34]
  assign _T_1894 = ab2_1_6 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2198 = _T_1894 ? 16'hcc : ab2_1_6; // @[loaf.scala 298:37]
  assign _T_1896 = macs_1_6_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_1898 = BFbuf_e > AEbuf_2_6_e; // @[loaf.scala 292:22]
  assign _T_1900 = AEbuf_2_6_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_1902 = AEbuf_2_6_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_1904 = BFbuf_a - AEbuf_2_6_a; // @[loaf.scala 295:34]
  assign _T_1906 = ab2_2_6 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2201 = _T_1906 ? 16'hcc : ab2_2_6; // @[loaf.scala 298:37]
  assign _T_1908 = macs_2_6_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_1910 = BFbuf_e > AEbuf_3_6_e; // @[loaf.scala 292:22]
  assign _T_1912 = AEbuf_3_6_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_1914 = AEbuf_3_6_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_1916 = BFbuf_a - AEbuf_3_6_a; // @[loaf.scala 295:34]
  assign _T_1918 = ab2_3_6 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2204 = _T_1918 ? 16'hcc : ab2_3_6; // @[loaf.scala 298:37]
  assign _T_1920 = macs_3_6_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_1922 = BFbuf_e > AEbuf_4_6_e; // @[loaf.scala 292:22]
  assign _T_1924 = AEbuf_4_6_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_1926 = AEbuf_4_6_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_1928 = BFbuf_a - AEbuf_4_6_a; // @[loaf.scala 295:34]
  assign _T_1930 = ab2_4_6 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2207 = _T_1930 ? 16'hcc : ab2_4_6; // @[loaf.scala 298:37]
  assign _T_1932 = macs_4_6_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_1934 = BFbuf_e > AEbuf_5_6_e; // @[loaf.scala 292:22]
  assign _T_1936 = AEbuf_5_6_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_1938 = AEbuf_5_6_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_1940 = BFbuf_a - AEbuf_5_6_a; // @[loaf.scala 295:34]
  assign _T_1942 = ab2_5_6 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2210 = _T_1942 ? 16'hcc : ab2_5_6; // @[loaf.scala 298:37]
  assign _T_1944 = macs_5_6_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_1946 = BFbuf_e > AEbuf_6_6_e; // @[loaf.scala 292:22]
  assign _T_1948 = AEbuf_6_6_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_1950 = AEbuf_6_6_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_1952 = BFbuf_a - AEbuf_6_6_a; // @[loaf.scala 295:34]
  assign _T_1954 = ab2_6_6 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2213 = _T_1954 ? 16'hcc : ab2_6_6; // @[loaf.scala 298:37]
  assign _T_1956 = macs_6_6_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_1958 = BFbuf_e > AEbuf_7_6_e; // @[loaf.scala 292:22]
  assign _T_1960 = AEbuf_7_6_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_1962 = AEbuf_7_6_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_1964 = BFbuf_a - AEbuf_7_6_a; // @[loaf.scala 295:34]
  assign _T_1966 = ab2_7_6 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2216 = _T_1966 ? 16'hcc : ab2_7_6; // @[loaf.scala 298:37]
  assign _T_1968 = macs_7_6_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_1970 = $signed(_T_1884) < $signed(_T_1896); // @[loaf.scala 327:24]
  assign _GEN_2217 = _T_1970 ? $signed(_T_1884) : $signed(_T_1896); // @[loaf.scala 327:29]
  assign _T_1972 = $signed(_T_1908) < $signed(_T_1920); // @[loaf.scala 327:24]
  assign _GEN_2218 = _T_1972 ? $signed(_T_1908) : $signed(_T_1920); // @[loaf.scala 327:29]
  assign _T_1974 = $signed(_T_1932) < $signed(_T_1944); // @[loaf.scala 327:24]
  assign _GEN_2219 = _T_1974 ? $signed(_T_1932) : $signed(_T_1944); // @[loaf.scala 327:29]
  assign _T_1976 = $signed(_T_1956) < $signed(_T_1968); // @[loaf.scala 327:24]
  assign _GEN_2220 = _T_1976 ? $signed(_T_1956) : $signed(_T_1968); // @[loaf.scala 327:29]
  assign _T_1978 = $signed(tm8_0_6) < $signed(tm8_1_6); // @[loaf.scala 327:24]
  assign _T_1980 = $signed(tm8_2_6) < $signed(tm8_3_6); // @[loaf.scala 327:24]
  assign _T_1982 = $signed(tm9_0_6) < $signed(tm9_1_6); // @[loaf.scala 327:24]
  assign _T_1984 = $signed(tmc_0_6) < $signed(best_6); // @[loaf.scala 354:43]
  assign _T_1985 = _T_448 | _T_1984; // @[loaf.scala 354:35]
  assign _T_1987 = BFbuf_e > AEbuf_0_7_e; // @[loaf.scala 292:22]
  assign _T_1989 = AEbuf_0_7_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_1991 = AEbuf_0_7_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_1993 = BFbuf_a - AEbuf_0_7_a; // @[loaf.scala 295:34]
  assign _T_1995 = ab2_0_7 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2227 = _T_1995 ? 16'hcc : ab2_0_7; // @[loaf.scala 298:37]
  assign _T_1997 = macs_0_7_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_1999 = BFbuf_e > AEbuf_1_7_e; // @[loaf.scala 292:22]
  assign _T_2001 = AEbuf_1_7_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_2003 = AEbuf_1_7_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_2005 = BFbuf_a - AEbuf_1_7_a; // @[loaf.scala 295:34]
  assign _T_2007 = ab2_1_7 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2230 = _T_2007 ? 16'hcc : ab2_1_7; // @[loaf.scala 298:37]
  assign _T_2009 = macs_1_7_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_2011 = BFbuf_e > AEbuf_2_7_e; // @[loaf.scala 292:22]
  assign _T_2013 = AEbuf_2_7_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_2015 = AEbuf_2_7_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_2017 = BFbuf_a - AEbuf_2_7_a; // @[loaf.scala 295:34]
  assign _T_2019 = ab2_2_7 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2233 = _T_2019 ? 16'hcc : ab2_2_7; // @[loaf.scala 298:37]
  assign _T_2021 = macs_2_7_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_2023 = BFbuf_e > AEbuf_3_7_e; // @[loaf.scala 292:22]
  assign _T_2025 = AEbuf_3_7_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_2027 = AEbuf_3_7_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_2029 = BFbuf_a - AEbuf_3_7_a; // @[loaf.scala 295:34]
  assign _T_2031 = ab2_3_7 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2236 = _T_2031 ? 16'hcc : ab2_3_7; // @[loaf.scala 298:37]
  assign _T_2033 = macs_3_7_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_2035 = BFbuf_e > AEbuf_4_7_e; // @[loaf.scala 292:22]
  assign _T_2037 = AEbuf_4_7_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_2039 = AEbuf_4_7_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_2041 = BFbuf_a - AEbuf_4_7_a; // @[loaf.scala 295:34]
  assign _T_2043 = ab2_4_7 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2239 = _T_2043 ? 16'hcc : ab2_4_7; // @[loaf.scala 298:37]
  assign _T_2045 = macs_4_7_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_2047 = BFbuf_e > AEbuf_5_7_e; // @[loaf.scala 292:22]
  assign _T_2049 = AEbuf_5_7_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_2051 = AEbuf_5_7_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_2053 = BFbuf_a - AEbuf_5_7_a; // @[loaf.scala 295:34]
  assign _T_2055 = ab2_5_7 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2242 = _T_2055 ? 16'hcc : ab2_5_7; // @[loaf.scala 298:37]
  assign _T_2057 = macs_5_7_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_2059 = BFbuf_e > AEbuf_6_7_e; // @[loaf.scala 292:22]
  assign _T_2061 = AEbuf_6_7_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_2063 = AEbuf_6_7_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_2065 = BFbuf_a - AEbuf_6_7_a; // @[loaf.scala 295:34]
  assign _T_2067 = ab2_6_7 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2245 = _T_2067 ? 16'hcc : ab2_6_7; // @[loaf.scala 298:37]
  assign _T_2069 = macs_6_7_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_2071 = BFbuf_e > AEbuf_7_7_e; // @[loaf.scala 292:22]
  assign _T_2073 = AEbuf_7_7_a - BFbuf_a; // @[loaf.scala 294:33]
  assign _T_2075 = AEbuf_7_7_a < BFbuf_a; // @[loaf.scala 295:21]
  assign _T_2077 = BFbuf_a - AEbuf_7_7_a; // @[loaf.scala 295:34]
  assign _T_2079 = ab2_7_7 > 16'hcc; // @[loaf.scala 298:29]
  assign _GEN_2248 = _T_2079 ? 16'hcc : ab2_7_7; // @[loaf.scala 298:37]
  assign _T_2081 = macs_7_7_io_r[31:10]; // @[loaf.scala 316:29]
  assign _T_2083 = $signed(_T_1997) < $signed(_T_2009); // @[loaf.scala 327:24]
  assign _GEN_2249 = _T_2083 ? $signed(_T_1997) : $signed(_T_2009); // @[loaf.scala 327:29]
  assign _T_2085 = $signed(_T_2021) < $signed(_T_2033); // @[loaf.scala 327:24]
  assign _GEN_2250 = _T_2085 ? $signed(_T_2021) : $signed(_T_2033); // @[loaf.scala 327:29]
  assign _T_2087 = $signed(_T_2045) < $signed(_T_2057); // @[loaf.scala 327:24]
  assign _GEN_2251 = _T_2087 ? $signed(_T_2045) : $signed(_T_2057); // @[loaf.scala 327:29]
  assign _T_2089 = $signed(_T_2069) < $signed(_T_2081); // @[loaf.scala 327:24]
  assign _GEN_2252 = _T_2089 ? $signed(_T_2069) : $signed(_T_2081); // @[loaf.scala 327:29]
  assign _T_2091 = $signed(tm8_0_7) < $signed(tm8_1_7); // @[loaf.scala 327:24]
  assign _T_2093 = $signed(tm8_2_7) < $signed(tm8_3_7); // @[loaf.scala 327:24]
  assign _T_2095 = $signed(tm9_0_7) < $signed(tm9_1_7); // @[loaf.scala 327:24]
  assign _T_2097 = $signed(tmc_0_7) < $signed(best_7); // @[loaf.scala 354:43]
  assign _T_2098 = _T_448 | _T_2097; // @[loaf.scala 354:35]
  assign _T_2102 = r != 2'h2; // @[loaf.scala 363:20]
  assign _T_2104 = r + 2'h1; // @[loaf.scala 364:20]
  assign _T_2105 = c != 2'h2; // @[loaf.scala 367:22]
  assign _T_2107 = c + 2'h1; // @[loaf.scala 368:22]
  assign _T_2108 = islice != 9'h113; // @[loaf.scala 375:31]
  assign _T_2110 = islice + 9'h1; // @[loaf.scala 376:36]
  assign _T_2112 = _T_405 == 1'h0; // @[loaf.scala 388:75]
  assign _T_2114 = _T_406 == 1'h0; // @[loaf.scala 388:75]
  assign _T_2115 = _T_2112 & _T_2114; // @[loaf.scala 388:72]
  assign _T_2116 = _T_407 == 1'h0; // @[loaf.scala 388:75]
  assign _T_2117 = _T_2115 & _T_2116; // @[loaf.scala 388:72]
  assign _T_2118 = _T_408 == 1'h0; // @[loaf.scala 388:75]
  assign _T_2119 = _T_2117 & _T_2118; // @[loaf.scala 388:72]
  assign _T_2120 = _T_409 == 1'h0; // @[loaf.scala 388:75]
  assign _T_2121 = _T_2119 & _T_2120; // @[loaf.scala 388:72]
  assign _T_2122 = _T_410 == 1'h0; // @[loaf.scala 388:75]
  assign _T_2123 = _T_2121 & _T_2122; // @[loaf.scala 388:72]
  assign _T_2124 = _T_411 == 1'h0; // @[loaf.scala 388:75]
  assign _T_2125 = _T_2123 & _T_2124; // @[loaf.scala 388:72]
  assign _T_2126 = _T_412 == 1'h0; // @[loaf.scala 388:75]
  assign _T_2127 = _T_2125 & _T_2126; // @[loaf.scala 388:72]
  assign _T_2128 = _T_413 == 1'h0; // @[loaf.scala 388:75]
  assign _T_2129 = _T_2127 & _T_2128; // @[loaf.scala 388:72]
  assign _T_2130 = _T_414 == 1'h0; // @[loaf.scala 388:75]
  assign _T_2131 = _T_2129 & _T_2130; // @[loaf.scala 388:72]
  assign _T_2132 = _T_415 == 1'h0; // @[loaf.scala 388:75]
  assign _T_2133 = _T_2131 & _T_2132; // @[loaf.scala 388:72]
  assign _T_2134 = _T_416 == 1'h0; // @[loaf.scala 388:75]
  assign _T_2135 = _T_2133 & _T_2134; // @[loaf.scala 388:72]
  assign _T_2136 = _T_417 == 1'h0; // @[loaf.scala 388:75]
  assign _T_2137 = _T_2135 & _T_2136; // @[loaf.scala 388:72]
  assign _T_2138 = _T_418 == 1'h0; // @[loaf.scala 388:75]
  assign _T_2139 = _T_2137 & _T_2138; // @[loaf.scala 388:72]
  assign _GEN_2323 = _T_463 ? _T_434 : 1'h0; // @[loaf.scala 246:49]
  assign _GEN_2324 = _T_463 ? _GEN_1763 : 1'h0; // @[loaf.scala 246:49]
  assign _GEN_2365 = _T_463 ? _T_487 : 1'h0; // @[loaf.scala 246:49]
  assign _GEN_2370 = _T_463 ? _T_466 : 1'h0; // @[loaf.scala 246:49]
  assign _GEN_2573 = _T_463 ? $signed(_T_1205) : $signed(26'sh0); // @[loaf.scala 246:49]
  assign _GEN_2574 = _T_463 ? mx2_0_0 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2575 = _T_463 ? _GEN_2003 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2578 = _T_463 ? $signed(_T_1217) : $signed(26'sh0); // @[loaf.scala 246:49]
  assign _GEN_2579 = _T_463 ? mx2_1_0 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2580 = _T_463 ? _GEN_2006 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2583 = _T_463 ? $signed(_T_1229) : $signed(26'sh0); // @[loaf.scala 246:49]
  assign _GEN_2584 = _T_463 ? mx2_2_0 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2585 = _T_463 ? _GEN_2009 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2588 = _T_463 ? $signed(_T_1241) : $signed(26'sh0); // @[loaf.scala 246:49]
  assign _GEN_2589 = _T_463 ? mx2_3_0 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2590 = _T_463 ? _GEN_2012 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2593 = _T_463 ? $signed(_T_1253) : $signed(26'sh0); // @[loaf.scala 246:49]
  assign _GEN_2594 = _T_463 ? mx2_4_0 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2595 = _T_463 ? _GEN_2015 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2598 = _T_463 ? $signed(_T_1265) : $signed(26'sh0); // @[loaf.scala 246:49]
  assign _GEN_2599 = _T_463 ? mx2_5_0 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2600 = _T_463 ? _GEN_2018 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2603 = _T_463 ? $signed(_T_1277) : $signed(26'sh0); // @[loaf.scala 246:49]
  assign _GEN_2604 = _T_463 ? mx2_6_0 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2605 = _T_463 ? _GEN_2021 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2608 = _T_463 ? $signed(_T_1289) : $signed(26'sh0); // @[loaf.scala 246:49]
  assign _GEN_2609 = _T_463 ? mx2_7_0 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2610 = _T_463 ? _GEN_2024 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2611 = _T_463 ? $signed(_GEN_2025) : $signed({{6{tm8_0_0[15]}},tm8_0_0}); // @[loaf.scala 246:49]
  assign _GEN_2612 = _T_463 ? $signed(_GEN_2026) : $signed({{6{tm8_1_0[15]}},tm8_1_0}); // @[loaf.scala 246:49]
  assign _GEN_2613 = _T_463 ? $signed(_GEN_2027) : $signed({{6{tm8_2_0[15]}},tm8_2_0}); // @[loaf.scala 246:49]
  assign _GEN_2614 = _T_463 ? $signed(_GEN_2028) : $signed({{6{tm8_3_0[15]}},tm8_3_0}); // @[loaf.scala 246:49]
  assign _GEN_2624 = _T_463 ? mx2_0_1 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2625 = _T_463 ? _GEN_2035 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2629 = _T_463 ? mx2_1_1 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2630 = _T_463 ? _GEN_2038 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2634 = _T_463 ? mx2_2_1 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2635 = _T_463 ? _GEN_2041 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2639 = _T_463 ? mx2_3_1 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2640 = _T_463 ? _GEN_2044 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2644 = _T_463 ? mx2_4_1 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2645 = _T_463 ? _GEN_2047 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2649 = _T_463 ? mx2_5_1 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2650 = _T_463 ? _GEN_2050 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2654 = _T_463 ? mx2_6_1 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2655 = _T_463 ? _GEN_2053 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2659 = _T_463 ? mx2_7_1 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2660 = _T_463 ? _GEN_2056 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2661 = _T_463 ? $signed(_GEN_2057) : $signed({{6{tm8_0_1[15]}},tm8_0_1}); // @[loaf.scala 246:49]
  assign _GEN_2662 = _T_463 ? $signed(_GEN_2058) : $signed({{6{tm8_1_1[15]}},tm8_1_1}); // @[loaf.scala 246:49]
  assign _GEN_2663 = _T_463 ? $signed(_GEN_2059) : $signed({{6{tm8_2_1[15]}},tm8_2_1}); // @[loaf.scala 246:49]
  assign _GEN_2664 = _T_463 ? $signed(_GEN_2060) : $signed({{6{tm8_3_1[15]}},tm8_3_1}); // @[loaf.scala 246:49]
  assign _GEN_2674 = _T_463 ? mx2_0_2 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2675 = _T_463 ? _GEN_2067 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2679 = _T_463 ? mx2_1_2 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2680 = _T_463 ? _GEN_2070 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2684 = _T_463 ? mx2_2_2 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2685 = _T_463 ? _GEN_2073 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2689 = _T_463 ? mx2_3_2 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2690 = _T_463 ? _GEN_2076 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2694 = _T_463 ? mx2_4_2 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2695 = _T_463 ? _GEN_2079 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2699 = _T_463 ? mx2_5_2 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2700 = _T_463 ? _GEN_2082 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2704 = _T_463 ? mx2_6_2 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2705 = _T_463 ? _GEN_2085 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2709 = _T_463 ? mx2_7_2 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2710 = _T_463 ? _GEN_2088 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2711 = _T_463 ? $signed(_GEN_2089) : $signed({{6{tm8_0_2[15]}},tm8_0_2}); // @[loaf.scala 246:49]
  assign _GEN_2712 = _T_463 ? $signed(_GEN_2090) : $signed({{6{tm8_1_2[15]}},tm8_1_2}); // @[loaf.scala 246:49]
  assign _GEN_2713 = _T_463 ? $signed(_GEN_2091) : $signed({{6{tm8_2_2[15]}},tm8_2_2}); // @[loaf.scala 246:49]
  assign _GEN_2714 = _T_463 ? $signed(_GEN_2092) : $signed({{6{tm8_3_2[15]}},tm8_3_2}); // @[loaf.scala 246:49]
  assign _GEN_2724 = _T_463 ? mx2_0_3 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2725 = _T_463 ? _GEN_2099 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2729 = _T_463 ? mx2_1_3 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2730 = _T_463 ? _GEN_2102 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2734 = _T_463 ? mx2_2_3 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2735 = _T_463 ? _GEN_2105 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2739 = _T_463 ? mx2_3_3 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2740 = _T_463 ? _GEN_2108 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2744 = _T_463 ? mx2_4_3 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2745 = _T_463 ? _GEN_2111 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2749 = _T_463 ? mx2_5_3 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2750 = _T_463 ? _GEN_2114 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2754 = _T_463 ? mx2_6_3 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2755 = _T_463 ? _GEN_2117 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2759 = _T_463 ? mx2_7_3 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2760 = _T_463 ? _GEN_2120 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2761 = _T_463 ? $signed(_GEN_2121) : $signed({{6{tm8_0_3[15]}},tm8_0_3}); // @[loaf.scala 246:49]
  assign _GEN_2762 = _T_463 ? $signed(_GEN_2122) : $signed({{6{tm8_1_3[15]}},tm8_1_3}); // @[loaf.scala 246:49]
  assign _GEN_2763 = _T_463 ? $signed(_GEN_2123) : $signed({{6{tm8_2_3[15]}},tm8_2_3}); // @[loaf.scala 246:49]
  assign _GEN_2764 = _T_463 ? $signed(_GEN_2124) : $signed({{6{tm8_3_3[15]}},tm8_3_3}); // @[loaf.scala 246:49]
  assign _GEN_2774 = _T_463 ? mx2_0_4 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2775 = _T_463 ? _GEN_2131 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2779 = _T_463 ? mx2_1_4 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2780 = _T_463 ? _GEN_2134 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2784 = _T_463 ? mx2_2_4 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2785 = _T_463 ? _GEN_2137 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2789 = _T_463 ? mx2_3_4 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2790 = _T_463 ? _GEN_2140 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2794 = _T_463 ? mx2_4_4 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2795 = _T_463 ? _GEN_2143 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2799 = _T_463 ? mx2_5_4 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2800 = _T_463 ? _GEN_2146 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2804 = _T_463 ? mx2_6_4 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2805 = _T_463 ? _GEN_2149 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2809 = _T_463 ? mx2_7_4 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2810 = _T_463 ? _GEN_2152 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2811 = _T_463 ? $signed(_GEN_2153) : $signed({{6{tm8_0_4[15]}},tm8_0_4}); // @[loaf.scala 246:49]
  assign _GEN_2812 = _T_463 ? $signed(_GEN_2154) : $signed({{6{tm8_1_4[15]}},tm8_1_4}); // @[loaf.scala 246:49]
  assign _GEN_2813 = _T_463 ? $signed(_GEN_2155) : $signed({{6{tm8_2_4[15]}},tm8_2_4}); // @[loaf.scala 246:49]
  assign _GEN_2814 = _T_463 ? $signed(_GEN_2156) : $signed({{6{tm8_3_4[15]}},tm8_3_4}); // @[loaf.scala 246:49]
  assign _GEN_2824 = _T_463 ? mx2_0_5 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2825 = _T_463 ? _GEN_2163 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2829 = _T_463 ? mx2_1_5 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2830 = _T_463 ? _GEN_2166 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2834 = _T_463 ? mx2_2_5 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2835 = _T_463 ? _GEN_2169 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2839 = _T_463 ? mx2_3_5 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2840 = _T_463 ? _GEN_2172 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2844 = _T_463 ? mx2_4_5 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2845 = _T_463 ? _GEN_2175 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2849 = _T_463 ? mx2_5_5 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2850 = _T_463 ? _GEN_2178 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2854 = _T_463 ? mx2_6_5 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2855 = _T_463 ? _GEN_2181 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2859 = _T_463 ? mx2_7_5 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2860 = _T_463 ? _GEN_2184 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2861 = _T_463 ? $signed(_GEN_2185) : $signed({{6{tm8_0_5[15]}},tm8_0_5}); // @[loaf.scala 246:49]
  assign _GEN_2862 = _T_463 ? $signed(_GEN_2186) : $signed({{6{tm8_1_5[15]}},tm8_1_5}); // @[loaf.scala 246:49]
  assign _GEN_2863 = _T_463 ? $signed(_GEN_2187) : $signed({{6{tm8_2_5[15]}},tm8_2_5}); // @[loaf.scala 246:49]
  assign _GEN_2864 = _T_463 ? $signed(_GEN_2188) : $signed({{6{tm8_3_5[15]}},tm8_3_5}); // @[loaf.scala 246:49]
  assign _GEN_2874 = _T_463 ? mx2_0_6 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2875 = _T_463 ? _GEN_2195 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2879 = _T_463 ? mx2_1_6 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2880 = _T_463 ? _GEN_2198 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2884 = _T_463 ? mx2_2_6 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2885 = _T_463 ? _GEN_2201 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2889 = _T_463 ? mx2_3_6 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2890 = _T_463 ? _GEN_2204 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2894 = _T_463 ? mx2_4_6 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2895 = _T_463 ? _GEN_2207 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2899 = _T_463 ? mx2_5_6 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2900 = _T_463 ? _GEN_2210 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2904 = _T_463 ? mx2_6_6 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2905 = _T_463 ? _GEN_2213 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2909 = _T_463 ? mx2_7_6 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2910 = _T_463 ? _GEN_2216 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2911 = _T_463 ? $signed(_GEN_2217) : $signed({{6{tm8_0_6[15]}},tm8_0_6}); // @[loaf.scala 246:49]
  assign _GEN_2912 = _T_463 ? $signed(_GEN_2218) : $signed({{6{tm8_1_6[15]}},tm8_1_6}); // @[loaf.scala 246:49]
  assign _GEN_2913 = _T_463 ? $signed(_GEN_2219) : $signed({{6{tm8_2_6[15]}},tm8_2_6}); // @[loaf.scala 246:49]
  assign _GEN_2914 = _T_463 ? $signed(_GEN_2220) : $signed({{6{tm8_3_6[15]}},tm8_3_6}); // @[loaf.scala 246:49]
  assign _GEN_2924 = _T_463 ? mx2_0_7 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2925 = _T_463 ? _GEN_2227 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2929 = _T_463 ? mx2_1_7 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2930 = _T_463 ? _GEN_2230 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2934 = _T_463 ? mx2_2_7 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2935 = _T_463 ? _GEN_2233 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2939 = _T_463 ? mx2_3_7 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2940 = _T_463 ? _GEN_2236 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2944 = _T_463 ? mx2_4_7 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2945 = _T_463 ? _GEN_2239 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2949 = _T_463 ? mx2_5_7 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2950 = _T_463 ? _GEN_2242 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2954 = _T_463 ? mx2_6_7 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2955 = _T_463 ? _GEN_2245 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2959 = _T_463 ? mx2_7_7 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2960 = _T_463 ? _GEN_2248 : 16'h0; // @[loaf.scala 246:49]
  assign _GEN_2961 = _T_463 ? $signed(_GEN_2249) : $signed({{6{tm8_0_7[15]}},tm8_0_7}); // @[loaf.scala 246:49]
  assign _GEN_2962 = _T_463 ? $signed(_GEN_2250) : $signed({{6{tm8_1_7[15]}},tm8_1_7}); // @[loaf.scala 246:49]
  assign _GEN_2963 = _T_463 ? $signed(_GEN_2251) : $signed({{6{tm8_2_7[15]}},tm8_2_7}); // @[loaf.scala 246:49]
  assign _GEN_2964 = _T_463 ? $signed(_GEN_2252) : $signed({{6{tm8_3_7[15]}},tm8_3_7}); // @[loaf.scala 246:49]
  assign _GEN_3036 = _T_452 ? _GEN_2323 : 1'h0; // @[loaf.scala 236:43]
  assign _GEN_3037 = _T_452 ? _GEN_2324 : 1'h0; // @[loaf.scala 236:43]
  assign _GEN_3078 = _T_452 ? _GEN_2365 : 1'h0; // @[loaf.scala 236:43]
  assign _GEN_3083 = _T_452 ? _GEN_2370 : 1'h0; // @[loaf.scala 236:43]
  assign _GEN_3285 = _T_452 ? _T_463 : 1'h0; // @[loaf.scala 236:43]
  assign _GEN_3286 = _T_452 ? $signed(_GEN_2573) : $signed(26'sh0); // @[loaf.scala 236:43]
  assign _GEN_3287 = _T_452 ? _GEN_2574 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3288 = _T_452 ? _GEN_2575 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3291 = _T_452 ? $signed(_GEN_2578) : $signed(26'sh0); // @[loaf.scala 236:43]
  assign _GEN_3292 = _T_452 ? _GEN_2579 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3293 = _T_452 ? _GEN_2580 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3296 = _T_452 ? $signed(_GEN_2583) : $signed(26'sh0); // @[loaf.scala 236:43]
  assign _GEN_3297 = _T_452 ? _GEN_2584 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3298 = _T_452 ? _GEN_2585 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3301 = _T_452 ? $signed(_GEN_2588) : $signed(26'sh0); // @[loaf.scala 236:43]
  assign _GEN_3302 = _T_452 ? _GEN_2589 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3303 = _T_452 ? _GEN_2590 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3306 = _T_452 ? $signed(_GEN_2593) : $signed(26'sh0); // @[loaf.scala 236:43]
  assign _GEN_3307 = _T_452 ? _GEN_2594 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3308 = _T_452 ? _GEN_2595 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3311 = _T_452 ? $signed(_GEN_2598) : $signed(26'sh0); // @[loaf.scala 236:43]
  assign _GEN_3312 = _T_452 ? _GEN_2599 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3313 = _T_452 ? _GEN_2600 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3316 = _T_452 ? $signed(_GEN_2603) : $signed(26'sh0); // @[loaf.scala 236:43]
  assign _GEN_3317 = _T_452 ? _GEN_2604 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3318 = _T_452 ? _GEN_2605 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3321 = _T_452 ? $signed(_GEN_2608) : $signed(26'sh0); // @[loaf.scala 236:43]
  assign _GEN_3322 = _T_452 ? _GEN_2609 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3323 = _T_452 ? _GEN_2610 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3324 = _T_452 ? $signed(_GEN_2611) : $signed({{6{tm8_0_0[15]}},tm8_0_0}); // @[loaf.scala 236:43]
  assign _GEN_3325 = _T_452 ? $signed(_GEN_2612) : $signed({{6{tm8_1_0[15]}},tm8_1_0}); // @[loaf.scala 236:43]
  assign _GEN_3326 = _T_452 ? $signed(_GEN_2613) : $signed({{6{tm8_2_0[15]}},tm8_2_0}); // @[loaf.scala 236:43]
  assign _GEN_3327 = _T_452 ? $signed(_GEN_2614) : $signed({{6{tm8_3_0[15]}},tm8_3_0}); // @[loaf.scala 236:43]
  assign _GEN_3337 = _T_452 ? _GEN_2624 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3338 = _T_452 ? _GEN_2625 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3342 = _T_452 ? _GEN_2629 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3343 = _T_452 ? _GEN_2630 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3347 = _T_452 ? _GEN_2634 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3348 = _T_452 ? _GEN_2635 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3352 = _T_452 ? _GEN_2639 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3353 = _T_452 ? _GEN_2640 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3357 = _T_452 ? _GEN_2644 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3358 = _T_452 ? _GEN_2645 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3362 = _T_452 ? _GEN_2649 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3363 = _T_452 ? _GEN_2650 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3367 = _T_452 ? _GEN_2654 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3368 = _T_452 ? _GEN_2655 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3372 = _T_452 ? _GEN_2659 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3373 = _T_452 ? _GEN_2660 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3374 = _T_452 ? $signed(_GEN_2661) : $signed({{6{tm8_0_1[15]}},tm8_0_1}); // @[loaf.scala 236:43]
  assign _GEN_3375 = _T_452 ? $signed(_GEN_2662) : $signed({{6{tm8_1_1[15]}},tm8_1_1}); // @[loaf.scala 236:43]
  assign _GEN_3376 = _T_452 ? $signed(_GEN_2663) : $signed({{6{tm8_2_1[15]}},tm8_2_1}); // @[loaf.scala 236:43]
  assign _GEN_3377 = _T_452 ? $signed(_GEN_2664) : $signed({{6{tm8_3_1[15]}},tm8_3_1}); // @[loaf.scala 236:43]
  assign _GEN_3387 = _T_452 ? _GEN_2674 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3388 = _T_452 ? _GEN_2675 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3392 = _T_452 ? _GEN_2679 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3393 = _T_452 ? _GEN_2680 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3397 = _T_452 ? _GEN_2684 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3398 = _T_452 ? _GEN_2685 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3402 = _T_452 ? _GEN_2689 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3403 = _T_452 ? _GEN_2690 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3407 = _T_452 ? _GEN_2694 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3408 = _T_452 ? _GEN_2695 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3412 = _T_452 ? _GEN_2699 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3413 = _T_452 ? _GEN_2700 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3417 = _T_452 ? _GEN_2704 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3418 = _T_452 ? _GEN_2705 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3422 = _T_452 ? _GEN_2709 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3423 = _T_452 ? _GEN_2710 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3424 = _T_452 ? $signed(_GEN_2711) : $signed({{6{tm8_0_2[15]}},tm8_0_2}); // @[loaf.scala 236:43]
  assign _GEN_3425 = _T_452 ? $signed(_GEN_2712) : $signed({{6{tm8_1_2[15]}},tm8_1_2}); // @[loaf.scala 236:43]
  assign _GEN_3426 = _T_452 ? $signed(_GEN_2713) : $signed({{6{tm8_2_2[15]}},tm8_2_2}); // @[loaf.scala 236:43]
  assign _GEN_3427 = _T_452 ? $signed(_GEN_2714) : $signed({{6{tm8_3_2[15]}},tm8_3_2}); // @[loaf.scala 236:43]
  assign _GEN_3437 = _T_452 ? _GEN_2724 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3438 = _T_452 ? _GEN_2725 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3442 = _T_452 ? _GEN_2729 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3443 = _T_452 ? _GEN_2730 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3447 = _T_452 ? _GEN_2734 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3448 = _T_452 ? _GEN_2735 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3452 = _T_452 ? _GEN_2739 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3453 = _T_452 ? _GEN_2740 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3457 = _T_452 ? _GEN_2744 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3458 = _T_452 ? _GEN_2745 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3462 = _T_452 ? _GEN_2749 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3463 = _T_452 ? _GEN_2750 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3467 = _T_452 ? _GEN_2754 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3468 = _T_452 ? _GEN_2755 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3472 = _T_452 ? _GEN_2759 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3473 = _T_452 ? _GEN_2760 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3474 = _T_452 ? $signed(_GEN_2761) : $signed({{6{tm8_0_3[15]}},tm8_0_3}); // @[loaf.scala 236:43]
  assign _GEN_3475 = _T_452 ? $signed(_GEN_2762) : $signed({{6{tm8_1_3[15]}},tm8_1_3}); // @[loaf.scala 236:43]
  assign _GEN_3476 = _T_452 ? $signed(_GEN_2763) : $signed({{6{tm8_2_3[15]}},tm8_2_3}); // @[loaf.scala 236:43]
  assign _GEN_3477 = _T_452 ? $signed(_GEN_2764) : $signed({{6{tm8_3_3[15]}},tm8_3_3}); // @[loaf.scala 236:43]
  assign _GEN_3487 = _T_452 ? _GEN_2774 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3488 = _T_452 ? _GEN_2775 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3492 = _T_452 ? _GEN_2779 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3493 = _T_452 ? _GEN_2780 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3497 = _T_452 ? _GEN_2784 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3498 = _T_452 ? _GEN_2785 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3502 = _T_452 ? _GEN_2789 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3503 = _T_452 ? _GEN_2790 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3507 = _T_452 ? _GEN_2794 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3508 = _T_452 ? _GEN_2795 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3512 = _T_452 ? _GEN_2799 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3513 = _T_452 ? _GEN_2800 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3517 = _T_452 ? _GEN_2804 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3518 = _T_452 ? _GEN_2805 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3522 = _T_452 ? _GEN_2809 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3523 = _T_452 ? _GEN_2810 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3524 = _T_452 ? $signed(_GEN_2811) : $signed({{6{tm8_0_4[15]}},tm8_0_4}); // @[loaf.scala 236:43]
  assign _GEN_3525 = _T_452 ? $signed(_GEN_2812) : $signed({{6{tm8_1_4[15]}},tm8_1_4}); // @[loaf.scala 236:43]
  assign _GEN_3526 = _T_452 ? $signed(_GEN_2813) : $signed({{6{tm8_2_4[15]}},tm8_2_4}); // @[loaf.scala 236:43]
  assign _GEN_3527 = _T_452 ? $signed(_GEN_2814) : $signed({{6{tm8_3_4[15]}},tm8_3_4}); // @[loaf.scala 236:43]
  assign _GEN_3537 = _T_452 ? _GEN_2824 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3538 = _T_452 ? _GEN_2825 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3542 = _T_452 ? _GEN_2829 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3543 = _T_452 ? _GEN_2830 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3547 = _T_452 ? _GEN_2834 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3548 = _T_452 ? _GEN_2835 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3552 = _T_452 ? _GEN_2839 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3553 = _T_452 ? _GEN_2840 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3557 = _T_452 ? _GEN_2844 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3558 = _T_452 ? _GEN_2845 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3562 = _T_452 ? _GEN_2849 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3563 = _T_452 ? _GEN_2850 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3567 = _T_452 ? _GEN_2854 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3568 = _T_452 ? _GEN_2855 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3572 = _T_452 ? _GEN_2859 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3573 = _T_452 ? _GEN_2860 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3574 = _T_452 ? $signed(_GEN_2861) : $signed({{6{tm8_0_5[15]}},tm8_0_5}); // @[loaf.scala 236:43]
  assign _GEN_3575 = _T_452 ? $signed(_GEN_2862) : $signed({{6{tm8_1_5[15]}},tm8_1_5}); // @[loaf.scala 236:43]
  assign _GEN_3576 = _T_452 ? $signed(_GEN_2863) : $signed({{6{tm8_2_5[15]}},tm8_2_5}); // @[loaf.scala 236:43]
  assign _GEN_3577 = _T_452 ? $signed(_GEN_2864) : $signed({{6{tm8_3_5[15]}},tm8_3_5}); // @[loaf.scala 236:43]
  assign _GEN_3587 = _T_452 ? _GEN_2874 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3588 = _T_452 ? _GEN_2875 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3592 = _T_452 ? _GEN_2879 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3593 = _T_452 ? _GEN_2880 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3597 = _T_452 ? _GEN_2884 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3598 = _T_452 ? _GEN_2885 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3602 = _T_452 ? _GEN_2889 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3603 = _T_452 ? _GEN_2890 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3607 = _T_452 ? _GEN_2894 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3608 = _T_452 ? _GEN_2895 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3612 = _T_452 ? _GEN_2899 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3613 = _T_452 ? _GEN_2900 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3617 = _T_452 ? _GEN_2904 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3618 = _T_452 ? _GEN_2905 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3622 = _T_452 ? _GEN_2909 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3623 = _T_452 ? _GEN_2910 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3624 = _T_452 ? $signed(_GEN_2911) : $signed({{6{tm8_0_6[15]}},tm8_0_6}); // @[loaf.scala 236:43]
  assign _GEN_3625 = _T_452 ? $signed(_GEN_2912) : $signed({{6{tm8_1_6[15]}},tm8_1_6}); // @[loaf.scala 236:43]
  assign _GEN_3626 = _T_452 ? $signed(_GEN_2913) : $signed({{6{tm8_2_6[15]}},tm8_2_6}); // @[loaf.scala 236:43]
  assign _GEN_3627 = _T_452 ? $signed(_GEN_2914) : $signed({{6{tm8_3_6[15]}},tm8_3_6}); // @[loaf.scala 236:43]
  assign _GEN_3637 = _T_452 ? _GEN_2924 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3638 = _T_452 ? _GEN_2925 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3642 = _T_452 ? _GEN_2929 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3643 = _T_452 ? _GEN_2930 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3647 = _T_452 ? _GEN_2934 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3648 = _T_452 ? _GEN_2935 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3652 = _T_452 ? _GEN_2939 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3653 = _T_452 ? _GEN_2940 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3657 = _T_452 ? _GEN_2944 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3658 = _T_452 ? _GEN_2945 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3662 = _T_452 ? _GEN_2949 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3663 = _T_452 ? _GEN_2950 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3667 = _T_452 ? _GEN_2954 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3668 = _T_452 ? _GEN_2955 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3672 = _T_452 ? _GEN_2959 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3673 = _T_452 ? _GEN_2960 : 16'h0; // @[loaf.scala 236:43]
  assign _GEN_3674 = _T_452 ? $signed(_GEN_2961) : $signed({{6{tm8_0_7[15]}},tm8_0_7}); // @[loaf.scala 236:43]
  assign _GEN_3675 = _T_452 ? $signed(_GEN_2962) : $signed({{6{tm8_1_7[15]}},tm8_1_7}); // @[loaf.scala 236:43]
  assign _GEN_3676 = _T_452 ? $signed(_GEN_2963) : $signed({{6{tm8_2_7[15]}},tm8_2_7}); // @[loaf.scala 236:43]
  assign _GEN_3677 = _T_452 ? $signed(_GEN_2964) : $signed({{6{tm8_3_7[15]}},tm8_3_7}); // @[loaf.scala 236:43]
  assign _GEN_3998 = _T_451 ? $signed(_GEN_3286) : $signed(26'sh0); // @[loaf.scala 234:29]
  assign _GEN_4003 = _T_451 ? $signed(_GEN_3291) : $signed(26'sh0); // @[loaf.scala 234:29]
  assign _GEN_4008 = _T_451 ? $signed(_GEN_3296) : $signed(26'sh0); // @[loaf.scala 234:29]
  assign _GEN_4013 = _T_451 ? $signed(_GEN_3301) : $signed(26'sh0); // @[loaf.scala 234:29]
  assign _GEN_4018 = _T_451 ? $signed(_GEN_3306) : $signed(26'sh0); // @[loaf.scala 234:29]
  assign _GEN_4023 = _T_451 ? $signed(_GEN_3311) : $signed(26'sh0); // @[loaf.scala 234:29]
  assign _GEN_4028 = _T_451 ? $signed(_GEN_3316) : $signed(26'sh0); // @[loaf.scala 234:29]
  assign _GEN_4033 = _T_451 ? $signed(_GEN_3321) : $signed(26'sh0); // @[loaf.scala 234:29]
  assign _GEN_4036 = _T_451 ? $signed(_GEN_3324) : $signed({{6{tm8_0_0[15]}},tm8_0_0}); // @[loaf.scala 234:29]
  assign _GEN_4037 = _T_451 ? $signed(_GEN_3325) : $signed({{6{tm8_1_0[15]}},tm8_1_0}); // @[loaf.scala 234:29]
  assign _GEN_4038 = _T_451 ? $signed(_GEN_3326) : $signed({{6{tm8_2_0[15]}},tm8_2_0}); // @[loaf.scala 234:29]
  assign _GEN_4039 = _T_451 ? $signed(_GEN_3327) : $signed({{6{tm8_3_0[15]}},tm8_3_0}); // @[loaf.scala 234:29]
  assign _GEN_4086 = _T_451 ? $signed(_GEN_3374) : $signed({{6{tm8_0_1[15]}},tm8_0_1}); // @[loaf.scala 234:29]
  assign _GEN_4087 = _T_451 ? $signed(_GEN_3375) : $signed({{6{tm8_1_1[15]}},tm8_1_1}); // @[loaf.scala 234:29]
  assign _GEN_4088 = _T_451 ? $signed(_GEN_3376) : $signed({{6{tm8_2_1[15]}},tm8_2_1}); // @[loaf.scala 234:29]
  assign _GEN_4089 = _T_451 ? $signed(_GEN_3377) : $signed({{6{tm8_3_1[15]}},tm8_3_1}); // @[loaf.scala 234:29]
  assign _GEN_4136 = _T_451 ? $signed(_GEN_3424) : $signed({{6{tm8_0_2[15]}},tm8_0_2}); // @[loaf.scala 234:29]
  assign _GEN_4137 = _T_451 ? $signed(_GEN_3425) : $signed({{6{tm8_1_2[15]}},tm8_1_2}); // @[loaf.scala 234:29]
  assign _GEN_4138 = _T_451 ? $signed(_GEN_3426) : $signed({{6{tm8_2_2[15]}},tm8_2_2}); // @[loaf.scala 234:29]
  assign _GEN_4139 = _T_451 ? $signed(_GEN_3427) : $signed({{6{tm8_3_2[15]}},tm8_3_2}); // @[loaf.scala 234:29]
  assign _GEN_4186 = _T_451 ? $signed(_GEN_3474) : $signed({{6{tm8_0_3[15]}},tm8_0_3}); // @[loaf.scala 234:29]
  assign _GEN_4187 = _T_451 ? $signed(_GEN_3475) : $signed({{6{tm8_1_3[15]}},tm8_1_3}); // @[loaf.scala 234:29]
  assign _GEN_4188 = _T_451 ? $signed(_GEN_3476) : $signed({{6{tm8_2_3[15]}},tm8_2_3}); // @[loaf.scala 234:29]
  assign _GEN_4189 = _T_451 ? $signed(_GEN_3477) : $signed({{6{tm8_3_3[15]}},tm8_3_3}); // @[loaf.scala 234:29]
  assign _GEN_4236 = _T_451 ? $signed(_GEN_3524) : $signed({{6{tm8_0_4[15]}},tm8_0_4}); // @[loaf.scala 234:29]
  assign _GEN_4237 = _T_451 ? $signed(_GEN_3525) : $signed({{6{tm8_1_4[15]}},tm8_1_4}); // @[loaf.scala 234:29]
  assign _GEN_4238 = _T_451 ? $signed(_GEN_3526) : $signed({{6{tm8_2_4[15]}},tm8_2_4}); // @[loaf.scala 234:29]
  assign _GEN_4239 = _T_451 ? $signed(_GEN_3527) : $signed({{6{tm8_3_4[15]}},tm8_3_4}); // @[loaf.scala 234:29]
  assign _GEN_4286 = _T_451 ? $signed(_GEN_3574) : $signed({{6{tm8_0_5[15]}},tm8_0_5}); // @[loaf.scala 234:29]
  assign _GEN_4287 = _T_451 ? $signed(_GEN_3575) : $signed({{6{tm8_1_5[15]}},tm8_1_5}); // @[loaf.scala 234:29]
  assign _GEN_4288 = _T_451 ? $signed(_GEN_3576) : $signed({{6{tm8_2_5[15]}},tm8_2_5}); // @[loaf.scala 234:29]
  assign _GEN_4289 = _T_451 ? $signed(_GEN_3577) : $signed({{6{tm8_3_5[15]}},tm8_3_5}); // @[loaf.scala 234:29]
  assign _GEN_4336 = _T_451 ? $signed(_GEN_3624) : $signed({{6{tm8_0_6[15]}},tm8_0_6}); // @[loaf.scala 234:29]
  assign _GEN_4337 = _T_451 ? $signed(_GEN_3625) : $signed({{6{tm8_1_6[15]}},tm8_1_6}); // @[loaf.scala 234:29]
  assign _GEN_4338 = _T_451 ? $signed(_GEN_3626) : $signed({{6{tm8_2_6[15]}},tm8_2_6}); // @[loaf.scala 234:29]
  assign _GEN_4339 = _T_451 ? $signed(_GEN_3627) : $signed({{6{tm8_3_6[15]}},tm8_3_6}); // @[loaf.scala 234:29]
  assign _GEN_4386 = _T_451 ? $signed(_GEN_3674) : $signed({{6{tm8_0_7[15]}},tm8_0_7}); // @[loaf.scala 234:29]
  assign _GEN_4387 = _T_451 ? $signed(_GEN_3675) : $signed({{6{tm8_1_7[15]}},tm8_1_7}); // @[loaf.scala 234:29]
  assign _GEN_4388 = _T_451 ? $signed(_GEN_3676) : $signed({{6{tm8_2_7[15]}},tm8_2_7}); // @[loaf.scala 234:29]
  assign _GEN_4389 = _T_451 ? $signed(_GEN_3677) : $signed({{6{tm8_3_7[15]}},tm8_3_7}); // @[loaf.scala 234:29]
  assign io_doneLoading = doneLoading; // @[loaf.scala 150:18]
  assign io_off_ready = _T_451 ? _GEN_3037 : 1'h0; // @[Decoupled.scala 69:20 loaf.scala 259:26]
  assign io_out_valid = _T_451 ? _GEN_3036 : 1'h0; // @[Decoupled.scala 53:20 loaf.scala 254:24]
  assign io_out_bits_0 = bestBufe_0; // @[loaf.scala 253:23]
  assign io_out_bits_1 = bestBufe_1; // @[loaf.scala 253:23]
  assign io_out_bits_2 = bestBufe_2; // @[loaf.scala 253:23]
  assign io_out_bits_3 = bestBufe_3; // @[loaf.scala 253:23]
  assign io_out_bits_4 = bestBufe_4; // @[loaf.scala 253:23]
  assign io_out_bits_5 = bestBufe_5; // @[loaf.scala 253:23]
  assign io_out_bits_6 = bestBufe_6; // @[loaf.scala 253:23]
  assign io_out_bits_7 = bestBufe_7; // @[loaf.scala 253:23]
  assign io_slc_ready = _T_2 ? _GEN_1309 : 1'h0; // @[Decoupled.scala 69:20 loaf.scala 189:24]
  assign io_lof_ready = _T_451 ? _GEN_3078 : 1'h0; // @[Decoupled.scala 69:20 loaf.scala 268:24]
  assign macs_0_0_clock = clock;
  assign macs_0_0_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_0_0_io_a = _T_451 ? _GEN_3287 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_0_0_io_b = _T_451 ? _GEN_3288 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_0_0_io_o = {{6{_GEN_3998[25]}},_GEN_3998}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign macs_0_1_clock = clock;
  assign macs_0_1_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_0_1_io_a = _T_451 ? _GEN_3337 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_0_1_io_b = _T_451 ? _GEN_3338 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_0_1_io_o = {{6{_GEN_3998[25]}},_GEN_3998}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign macs_0_2_clock = clock;
  assign macs_0_2_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_0_2_io_a = _T_451 ? _GEN_3387 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_0_2_io_b = _T_451 ? _GEN_3388 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_0_2_io_o = {{6{_GEN_3998[25]}},_GEN_3998}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign macs_0_3_clock = clock;
  assign macs_0_3_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_0_3_io_a = _T_451 ? _GEN_3437 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_0_3_io_b = _T_451 ? _GEN_3438 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_0_3_io_o = {{6{_GEN_3998[25]}},_GEN_3998}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign macs_0_4_clock = clock;
  assign macs_0_4_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_0_4_io_a = _T_451 ? _GEN_3487 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_0_4_io_b = _T_451 ? _GEN_3488 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_0_4_io_o = {{6{_GEN_3998[25]}},_GEN_3998}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign macs_0_5_clock = clock;
  assign macs_0_5_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_0_5_io_a = _T_451 ? _GEN_3537 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_0_5_io_b = _T_451 ? _GEN_3538 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_0_5_io_o = {{6{_GEN_3998[25]}},_GEN_3998}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign macs_0_6_clock = clock;
  assign macs_0_6_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_0_6_io_a = _T_451 ? _GEN_3587 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_0_6_io_b = _T_451 ? _GEN_3588 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_0_6_io_o = {{6{_GEN_3998[25]}},_GEN_3998}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign macs_0_7_clock = clock;
  assign macs_0_7_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_0_7_io_a = _T_451 ? _GEN_3637 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_0_7_io_b = _T_451 ? _GEN_3638 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_0_7_io_o = {{6{_GEN_3998[25]}},_GEN_3998}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign macs_1_0_clock = clock;
  assign macs_1_0_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_1_0_io_a = _T_451 ? _GEN_3292 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_1_0_io_b = _T_451 ? _GEN_3293 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_1_0_io_o = {{6{_GEN_4003[25]}},_GEN_4003}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign macs_1_1_clock = clock;
  assign macs_1_1_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_1_1_io_a = _T_451 ? _GEN_3342 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_1_1_io_b = _T_451 ? _GEN_3343 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_1_1_io_o = {{6{_GEN_4003[25]}},_GEN_4003}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign macs_1_2_clock = clock;
  assign macs_1_2_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_1_2_io_a = _T_451 ? _GEN_3392 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_1_2_io_b = _T_451 ? _GEN_3393 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_1_2_io_o = {{6{_GEN_4003[25]}},_GEN_4003}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign macs_1_3_clock = clock;
  assign macs_1_3_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_1_3_io_a = _T_451 ? _GEN_3442 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_1_3_io_b = _T_451 ? _GEN_3443 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_1_3_io_o = {{6{_GEN_4003[25]}},_GEN_4003}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign macs_1_4_clock = clock;
  assign macs_1_4_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_1_4_io_a = _T_451 ? _GEN_3492 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_1_4_io_b = _T_451 ? _GEN_3493 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_1_4_io_o = {{6{_GEN_4003[25]}},_GEN_4003}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign macs_1_5_clock = clock;
  assign macs_1_5_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_1_5_io_a = _T_451 ? _GEN_3542 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_1_5_io_b = _T_451 ? _GEN_3543 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_1_5_io_o = {{6{_GEN_4003[25]}},_GEN_4003}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign macs_1_6_clock = clock;
  assign macs_1_6_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_1_6_io_a = _T_451 ? _GEN_3592 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_1_6_io_b = _T_451 ? _GEN_3593 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_1_6_io_o = {{6{_GEN_4003[25]}},_GEN_4003}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign macs_1_7_clock = clock;
  assign macs_1_7_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_1_7_io_a = _T_451 ? _GEN_3642 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_1_7_io_b = _T_451 ? _GEN_3643 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_1_7_io_o = {{6{_GEN_4003[25]}},_GEN_4003}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign macs_2_0_clock = clock;
  assign macs_2_0_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_2_0_io_a = _T_451 ? _GEN_3297 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_2_0_io_b = _T_451 ? _GEN_3298 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_2_0_io_o = {{6{_GEN_4008[25]}},_GEN_4008}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign macs_2_1_clock = clock;
  assign macs_2_1_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_2_1_io_a = _T_451 ? _GEN_3347 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_2_1_io_b = _T_451 ? _GEN_3348 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_2_1_io_o = {{6{_GEN_4008[25]}},_GEN_4008}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign macs_2_2_clock = clock;
  assign macs_2_2_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_2_2_io_a = _T_451 ? _GEN_3397 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_2_2_io_b = _T_451 ? _GEN_3398 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_2_2_io_o = {{6{_GEN_4008[25]}},_GEN_4008}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign macs_2_3_clock = clock;
  assign macs_2_3_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_2_3_io_a = _T_451 ? _GEN_3447 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_2_3_io_b = _T_451 ? _GEN_3448 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_2_3_io_o = {{6{_GEN_4008[25]}},_GEN_4008}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign macs_2_4_clock = clock;
  assign macs_2_4_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_2_4_io_a = _T_451 ? _GEN_3497 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_2_4_io_b = _T_451 ? _GEN_3498 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_2_4_io_o = {{6{_GEN_4008[25]}},_GEN_4008}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign macs_2_5_clock = clock;
  assign macs_2_5_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_2_5_io_a = _T_451 ? _GEN_3547 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_2_5_io_b = _T_451 ? _GEN_3548 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_2_5_io_o = {{6{_GEN_4008[25]}},_GEN_4008}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign macs_2_6_clock = clock;
  assign macs_2_6_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_2_6_io_a = _T_451 ? _GEN_3597 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_2_6_io_b = _T_451 ? _GEN_3598 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_2_6_io_o = {{6{_GEN_4008[25]}},_GEN_4008}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign macs_2_7_clock = clock;
  assign macs_2_7_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_2_7_io_a = _T_451 ? _GEN_3647 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_2_7_io_b = _T_451 ? _GEN_3648 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_2_7_io_o = {{6{_GEN_4008[25]}},_GEN_4008}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign macs_3_0_clock = clock;
  assign macs_3_0_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_3_0_io_a = _T_451 ? _GEN_3302 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_3_0_io_b = _T_451 ? _GEN_3303 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_3_0_io_o = {{6{_GEN_4013[25]}},_GEN_4013}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign macs_3_1_clock = clock;
  assign macs_3_1_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_3_1_io_a = _T_451 ? _GEN_3352 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_3_1_io_b = _T_451 ? _GEN_3353 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_3_1_io_o = {{6{_GEN_4013[25]}},_GEN_4013}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign macs_3_2_clock = clock;
  assign macs_3_2_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_3_2_io_a = _T_451 ? _GEN_3402 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_3_2_io_b = _T_451 ? _GEN_3403 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_3_2_io_o = {{6{_GEN_4013[25]}},_GEN_4013}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign macs_3_3_clock = clock;
  assign macs_3_3_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_3_3_io_a = _T_451 ? _GEN_3452 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_3_3_io_b = _T_451 ? _GEN_3453 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_3_3_io_o = {{6{_GEN_4013[25]}},_GEN_4013}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign macs_3_4_clock = clock;
  assign macs_3_4_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_3_4_io_a = _T_451 ? _GEN_3502 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_3_4_io_b = _T_451 ? _GEN_3503 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_3_4_io_o = {{6{_GEN_4013[25]}},_GEN_4013}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign macs_3_5_clock = clock;
  assign macs_3_5_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_3_5_io_a = _T_451 ? _GEN_3552 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_3_5_io_b = _T_451 ? _GEN_3553 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_3_5_io_o = {{6{_GEN_4013[25]}},_GEN_4013}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign macs_3_6_clock = clock;
  assign macs_3_6_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_3_6_io_a = _T_451 ? _GEN_3602 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_3_6_io_b = _T_451 ? _GEN_3603 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_3_6_io_o = {{6{_GEN_4013[25]}},_GEN_4013}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign macs_3_7_clock = clock;
  assign macs_3_7_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_3_7_io_a = _T_451 ? _GEN_3652 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_3_7_io_b = _T_451 ? _GEN_3653 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_3_7_io_o = {{6{_GEN_4013[25]}},_GEN_4013}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign macs_4_0_clock = clock;
  assign macs_4_0_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_4_0_io_a = _T_451 ? _GEN_3307 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_4_0_io_b = _T_451 ? _GEN_3308 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_4_0_io_o = {{6{_GEN_4018[25]}},_GEN_4018}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign macs_4_1_clock = clock;
  assign macs_4_1_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_4_1_io_a = _T_451 ? _GEN_3357 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_4_1_io_b = _T_451 ? _GEN_3358 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_4_1_io_o = {{6{_GEN_4018[25]}},_GEN_4018}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign macs_4_2_clock = clock;
  assign macs_4_2_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_4_2_io_a = _T_451 ? _GEN_3407 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_4_2_io_b = _T_451 ? _GEN_3408 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_4_2_io_o = {{6{_GEN_4018[25]}},_GEN_4018}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign macs_4_3_clock = clock;
  assign macs_4_3_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_4_3_io_a = _T_451 ? _GEN_3457 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_4_3_io_b = _T_451 ? _GEN_3458 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_4_3_io_o = {{6{_GEN_4018[25]}},_GEN_4018}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign macs_4_4_clock = clock;
  assign macs_4_4_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_4_4_io_a = _T_451 ? _GEN_3507 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_4_4_io_b = _T_451 ? _GEN_3508 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_4_4_io_o = {{6{_GEN_4018[25]}},_GEN_4018}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign macs_4_5_clock = clock;
  assign macs_4_5_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_4_5_io_a = _T_451 ? _GEN_3557 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_4_5_io_b = _T_451 ? _GEN_3558 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_4_5_io_o = {{6{_GEN_4018[25]}},_GEN_4018}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign macs_4_6_clock = clock;
  assign macs_4_6_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_4_6_io_a = _T_451 ? _GEN_3607 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_4_6_io_b = _T_451 ? _GEN_3608 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_4_6_io_o = {{6{_GEN_4018[25]}},_GEN_4018}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign macs_4_7_clock = clock;
  assign macs_4_7_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_4_7_io_a = _T_451 ? _GEN_3657 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_4_7_io_b = _T_451 ? _GEN_3658 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_4_7_io_o = {{6{_GEN_4018[25]}},_GEN_4018}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign macs_5_0_clock = clock;
  assign macs_5_0_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_5_0_io_a = _T_451 ? _GEN_3312 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_5_0_io_b = _T_451 ? _GEN_3313 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_5_0_io_o = {{6{_GEN_4023[25]}},_GEN_4023}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign macs_5_1_clock = clock;
  assign macs_5_1_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_5_1_io_a = _T_451 ? _GEN_3362 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_5_1_io_b = _T_451 ? _GEN_3363 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_5_1_io_o = {{6{_GEN_4023[25]}},_GEN_4023}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign macs_5_2_clock = clock;
  assign macs_5_2_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_5_2_io_a = _T_451 ? _GEN_3412 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_5_2_io_b = _T_451 ? _GEN_3413 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_5_2_io_o = {{6{_GEN_4023[25]}},_GEN_4023}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign macs_5_3_clock = clock;
  assign macs_5_3_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_5_3_io_a = _T_451 ? _GEN_3462 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_5_3_io_b = _T_451 ? _GEN_3463 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_5_3_io_o = {{6{_GEN_4023[25]}},_GEN_4023}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign macs_5_4_clock = clock;
  assign macs_5_4_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_5_4_io_a = _T_451 ? _GEN_3512 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_5_4_io_b = _T_451 ? _GEN_3513 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_5_4_io_o = {{6{_GEN_4023[25]}},_GEN_4023}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign macs_5_5_clock = clock;
  assign macs_5_5_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_5_5_io_a = _T_451 ? _GEN_3562 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_5_5_io_b = _T_451 ? _GEN_3563 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_5_5_io_o = {{6{_GEN_4023[25]}},_GEN_4023}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign macs_5_6_clock = clock;
  assign macs_5_6_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_5_6_io_a = _T_451 ? _GEN_3612 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_5_6_io_b = _T_451 ? _GEN_3613 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_5_6_io_o = {{6{_GEN_4023[25]}},_GEN_4023}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign macs_5_7_clock = clock;
  assign macs_5_7_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_5_7_io_a = _T_451 ? _GEN_3662 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_5_7_io_b = _T_451 ? _GEN_3663 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_5_7_io_o = {{6{_GEN_4023[25]}},_GEN_4023}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign macs_6_0_clock = clock;
  assign macs_6_0_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_6_0_io_a = _T_451 ? _GEN_3317 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_6_0_io_b = _T_451 ? _GEN_3318 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_6_0_io_o = {{6{_GEN_4028[25]}},_GEN_4028}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign macs_6_1_clock = clock;
  assign macs_6_1_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_6_1_io_a = _T_451 ? _GEN_3367 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_6_1_io_b = _T_451 ? _GEN_3368 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_6_1_io_o = {{6{_GEN_4028[25]}},_GEN_4028}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign macs_6_2_clock = clock;
  assign macs_6_2_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_6_2_io_a = _T_451 ? _GEN_3417 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_6_2_io_b = _T_451 ? _GEN_3418 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_6_2_io_o = {{6{_GEN_4028[25]}},_GEN_4028}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign macs_6_3_clock = clock;
  assign macs_6_3_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_6_3_io_a = _T_451 ? _GEN_3467 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_6_3_io_b = _T_451 ? _GEN_3468 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_6_3_io_o = {{6{_GEN_4028[25]}},_GEN_4028}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign macs_6_4_clock = clock;
  assign macs_6_4_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_6_4_io_a = _T_451 ? _GEN_3517 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_6_4_io_b = _T_451 ? _GEN_3518 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_6_4_io_o = {{6{_GEN_4028[25]}},_GEN_4028}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign macs_6_5_clock = clock;
  assign macs_6_5_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_6_5_io_a = _T_451 ? _GEN_3567 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_6_5_io_b = _T_451 ? _GEN_3568 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_6_5_io_o = {{6{_GEN_4028[25]}},_GEN_4028}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign macs_6_6_clock = clock;
  assign macs_6_6_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_6_6_io_a = _T_451 ? _GEN_3617 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_6_6_io_b = _T_451 ? _GEN_3618 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_6_6_io_o = {{6{_GEN_4028[25]}},_GEN_4028}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign macs_6_7_clock = clock;
  assign macs_6_7_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_6_7_io_a = _T_451 ? _GEN_3667 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_6_7_io_b = _T_451 ? _GEN_3668 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_6_7_io_o = {{6{_GEN_4028[25]}},_GEN_4028}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign macs_7_0_clock = clock;
  assign macs_7_0_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_7_0_io_a = _T_451 ? _GEN_3322 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_7_0_io_b = _T_451 ? _GEN_3323 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_7_0_io_o = {{6{_GEN_4033[25]}},_GEN_4033}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign macs_7_1_clock = clock;
  assign macs_7_1_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_7_1_io_a = _T_451 ? _GEN_3372 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_7_1_io_b = _T_451 ? _GEN_3373 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_7_1_io_o = {{6{_GEN_4033[25]}},_GEN_4033}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign macs_7_2_clock = clock;
  assign macs_7_2_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_7_2_io_a = _T_451 ? _GEN_3422 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_7_2_io_b = _T_451 ? _GEN_3423 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_7_2_io_o = {{6{_GEN_4033[25]}},_GEN_4033}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign macs_7_3_clock = clock;
  assign macs_7_3_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_7_3_io_a = _T_451 ? _GEN_3472 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_7_3_io_b = _T_451 ? _GEN_3473 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_7_3_io_o = {{6{_GEN_4033[25]}},_GEN_4033}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign macs_7_4_clock = clock;
  assign macs_7_4_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_7_4_io_a = _T_451 ? _GEN_3522 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_7_4_io_b = _T_451 ? _GEN_3523 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_7_4_io_o = {{6{_GEN_4033[25]}},_GEN_4033}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign macs_7_5_clock = clock;
  assign macs_7_5_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_7_5_io_a = _T_451 ? _GEN_3572 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_7_5_io_b = _T_451 ? _GEN_3573 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_7_5_io_o = {{6{_GEN_4033[25]}},_GEN_4033}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign macs_7_6_clock = clock;
  assign macs_7_6_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_7_6_io_a = _T_451 ? _GEN_3622 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_7_6_io_b = _T_451 ? _GEN_3623 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_7_6_io_o = {{6{_GEN_4033[25]}},_GEN_4033}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign macs_7_7_clock = clock;
  assign macs_7_7_io_en = _T_451 ? _GEN_3285 : 1'h0; // @[loaf.scala 161:22 loaf.scala 300:30]
  assign macs_7_7_io_a = _T_451 ? _GEN_3672 : 16'h0; // @[loaf.scala 163:21 loaf.scala 303:29]
  assign macs_7_7_io_b = _T_451 ? _GEN_3673 : 16'h0; // @[loaf.scala 164:21 loaf.scala 304:29]
  assign macs_7_7_io_o = {{6{_GEN_4033[25]}},_GEN_4033}; // @[loaf.scala 165:21 loaf.scala 302:29]
  assign _GEN_4987 = _GEN_4036[15:0]; // @[loaf.scala 337:25]
  assign _GEN_4988 = _GEN_4086[15:0]; // @[loaf.scala 337:25]
  assign _GEN_4989 = _GEN_4136[15:0]; // @[loaf.scala 337:25]
  assign _GEN_4990 = _GEN_4186[15:0]; // @[loaf.scala 337:25]
  assign _GEN_4991 = _GEN_4236[15:0]; // @[loaf.scala 337:25]
  assign _GEN_4992 = _GEN_4286[15:0]; // @[loaf.scala 337:25]
  assign _GEN_4993 = _GEN_4336[15:0]; // @[loaf.scala 337:25]
  assign _GEN_4994 = _GEN_4386[15:0]; // @[loaf.scala 337:25]
  assign _GEN_4995 = _GEN_4037[15:0]; // @[loaf.scala 337:25]
  assign _GEN_4996 = _GEN_4087[15:0]; // @[loaf.scala 337:25]
  assign _GEN_4997 = _GEN_4137[15:0]; // @[loaf.scala 337:25]
  assign _GEN_4998 = _GEN_4187[15:0]; // @[loaf.scala 337:25]
  assign _GEN_4999 = _GEN_4237[15:0]; // @[loaf.scala 337:25]
  assign _GEN_5000 = _GEN_4287[15:0]; // @[loaf.scala 337:25]
  assign _GEN_5001 = _GEN_4337[15:0]; // @[loaf.scala 337:25]
  assign _GEN_5002 = _GEN_4387[15:0]; // @[loaf.scala 337:25]
  assign _GEN_5003 = _GEN_4038[15:0]; // @[loaf.scala 337:25]
  assign _GEN_5004 = _GEN_4088[15:0]; // @[loaf.scala 337:25]
  assign _GEN_5005 = _GEN_4138[15:0]; // @[loaf.scala 337:25]
  assign _GEN_5006 = _GEN_4188[15:0]; // @[loaf.scala 337:25]
  assign _GEN_5007 = _GEN_4238[15:0]; // @[loaf.scala 337:25]
  assign _GEN_5008 = _GEN_4288[15:0]; // @[loaf.scala 337:25]
  assign _GEN_5009 = _GEN_4338[15:0]; // @[loaf.scala 337:25]
  assign _GEN_5010 = _GEN_4388[15:0]; // @[loaf.scala 337:25]
  assign _GEN_5011 = _GEN_4039[15:0]; // @[loaf.scala 337:25]
  assign _GEN_5012 = _GEN_4089[15:0]; // @[loaf.scala 337:25]
  assign _GEN_5013 = _GEN_4139[15:0]; // @[loaf.scala 337:25]
  assign _GEN_5014 = _GEN_4189[15:0]; // @[loaf.scala 337:25]
  assign _GEN_5015 = _GEN_4239[15:0]; // @[loaf.scala 337:25]
  assign _GEN_5016 = _GEN_4289[15:0]; // @[loaf.scala 337:25]
  assign _GEN_5017 = _GEN_4339[15:0]; // @[loaf.scala 337:25]
  assign _GEN_5018 = _GEN_4389[15:0]; // @[loaf.scala 337:25]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_0_0[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_0_1[initvar] = _RAND_1[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_0_2[initvar] = _RAND_2[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_0_3[initvar] = _RAND_3[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_0_4[initvar] = _RAND_4[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_0_5[initvar] = _RAND_5[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_6 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_0_6[initvar] = _RAND_6[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_7 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_0_7[initvar] = _RAND_7[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_8 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_1_0[initvar] = _RAND_8[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_9 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_1_1[initvar] = _RAND_9[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_10 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_1_2[initvar] = _RAND_10[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_11 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_1_3[initvar] = _RAND_11[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_12 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_1_4[initvar] = _RAND_12[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_13 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_1_5[initvar] = _RAND_13[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_14 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_1_6[initvar] = _RAND_14[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_15 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_1_7[initvar] = _RAND_15[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_16 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_2_0[initvar] = _RAND_16[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_17 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_2_1[initvar] = _RAND_17[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_18 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_2_2[initvar] = _RAND_18[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_19 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_2_3[initvar] = _RAND_19[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_20 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_2_4[initvar] = _RAND_20[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_21 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_2_5[initvar] = _RAND_21[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_22 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_2_6[initvar] = _RAND_22[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_23 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_2_7[initvar] = _RAND_23[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_24 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_3_0[initvar] = _RAND_24[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_25 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_3_1[initvar] = _RAND_25[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_26 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_3_2[initvar] = _RAND_26[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_27 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_3_3[initvar] = _RAND_27[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_28 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_3_4[initvar] = _RAND_28[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_29 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_3_5[initvar] = _RAND_29[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_30 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_3_6[initvar] = _RAND_30[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_31 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_3_7[initvar] = _RAND_31[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_32 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_4_0[initvar] = _RAND_32[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_33 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_4_1[initvar] = _RAND_33[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_34 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_4_2[initvar] = _RAND_34[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_35 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_4_3[initvar] = _RAND_35[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_36 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_4_4[initvar] = _RAND_36[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_37 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_4_5[initvar] = _RAND_37[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_38 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_4_6[initvar] = _RAND_38[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_39 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_4_7[initvar] = _RAND_39[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_40 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_5_0[initvar] = _RAND_40[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_41 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_5_1[initvar] = _RAND_41[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_42 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_5_2[initvar] = _RAND_42[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_43 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_5_3[initvar] = _RAND_43[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_44 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_5_4[initvar] = _RAND_44[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_45 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_5_5[initvar] = _RAND_45[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_46 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_5_6[initvar] = _RAND_46[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_47 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_5_7[initvar] = _RAND_47[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_48 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_6_0[initvar] = _RAND_48[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_49 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_6_1[initvar] = _RAND_49[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_50 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_6_2[initvar] = _RAND_50[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_51 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_6_3[initvar] = _RAND_51[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_52 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_6_4[initvar] = _RAND_52[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_53 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_6_5[initvar] = _RAND_53[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_54 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_6_6[initvar] = _RAND_54[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_55 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_6_7[initvar] = _RAND_55[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_56 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_7_0[initvar] = _RAND_56[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_57 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_7_1[initvar] = _RAND_57[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_58 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_7_2[initvar] = _RAND_58[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_59 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_7_3[initvar] = _RAND_59[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_60 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_7_4[initvar] = _RAND_60[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_61 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_7_5[initvar] = _RAND_61[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_62 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_7_6[initvar] = _RAND_62[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_63 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    AE_7_7[initvar] = _RAND_63[31:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  islice = _RAND_64[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  done = _RAND_65[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  phase = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  offCLs_0_0 = _RAND_67[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  offCLs_0_1 = _RAND_68[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  offCLs_0_2 = _RAND_69[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  offCLs_0_3 = _RAND_70[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  offCLs_0_4 = _RAND_71[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  offCLs_0_5 = _RAND_72[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  offCLs_0_6 = _RAND_73[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  offCLs_0_7 = _RAND_74[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  offCLs_1_0 = _RAND_75[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  offCLs_1_1 = _RAND_76[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  offCLs_1_2 = _RAND_77[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  offCLs_1_3 = _RAND_78[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  offCLs_1_4 = _RAND_79[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  offCLs_1_5 = _RAND_80[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  offCLs_1_6 = _RAND_81[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  offCLs_1_7 = _RAND_82[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  offCLs_2_0 = _RAND_83[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  offCLs_2_1 = _RAND_84[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  offCLs_2_2 = _RAND_85[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  offCLs_2_3 = _RAND_86[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  offCLs_2_4 = _RAND_87[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  offCLs_2_5 = _RAND_88[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  offCLs_2_6 = _RAND_89[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  offCLs_2_7 = _RAND_90[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  offCLs_3_0 = _RAND_91[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  offCLs_3_1 = _RAND_92[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  offCLs_3_2 = _RAND_93[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  offCLs_3_3 = _RAND_94[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  offCLs_3_4 = _RAND_95[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  offCLs_3_5 = _RAND_96[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  offCLs_3_6 = _RAND_97[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  offCLs_3_7 = _RAND_98[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  o1_0 = _RAND_99[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  o1_1 = _RAND_100[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  o1_2 = _RAND_101[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  o1_3 = _RAND_102[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  o1_4 = _RAND_103[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  o1_5 = _RAND_104[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  o1_6 = _RAND_105[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  o1_7 = _RAND_106[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  o2_0 = _RAND_107[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  o2_1 = _RAND_108[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  o2_2 = _RAND_109[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  o2_3 = _RAND_110[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  o2_4 = _RAND_111[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  o2_5 = _RAND_112[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  o2_6 = _RAND_113[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  o2_7 = _RAND_114[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  mx2_0_0 = _RAND_115[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  mx2_0_1 = _RAND_116[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  mx2_0_2 = _RAND_117[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  mx2_0_3 = _RAND_118[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  mx2_0_4 = _RAND_119[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  mx2_0_5 = _RAND_120[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  mx2_0_6 = _RAND_121[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  mx2_0_7 = _RAND_122[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  mx2_1_0 = _RAND_123[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  mx2_1_1 = _RAND_124[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  mx2_1_2 = _RAND_125[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  mx2_1_3 = _RAND_126[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  mx2_1_4 = _RAND_127[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  mx2_1_5 = _RAND_128[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  mx2_1_6 = _RAND_129[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  mx2_1_7 = _RAND_130[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  mx2_2_0 = _RAND_131[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  mx2_2_1 = _RAND_132[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  mx2_2_2 = _RAND_133[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  mx2_2_3 = _RAND_134[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  mx2_2_4 = _RAND_135[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  mx2_2_5 = _RAND_136[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  mx2_2_6 = _RAND_137[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  mx2_2_7 = _RAND_138[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  mx2_3_0 = _RAND_139[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  mx2_3_1 = _RAND_140[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  mx2_3_2 = _RAND_141[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  mx2_3_3 = _RAND_142[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  mx2_3_4 = _RAND_143[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  mx2_3_5 = _RAND_144[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  mx2_3_6 = _RAND_145[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  mx2_3_7 = _RAND_146[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  mx2_4_0 = _RAND_147[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  mx2_4_1 = _RAND_148[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  mx2_4_2 = _RAND_149[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  mx2_4_3 = _RAND_150[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  mx2_4_4 = _RAND_151[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  mx2_4_5 = _RAND_152[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  mx2_4_6 = _RAND_153[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  mx2_4_7 = _RAND_154[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  mx2_5_0 = _RAND_155[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  mx2_5_1 = _RAND_156[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  mx2_5_2 = _RAND_157[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  mx2_5_3 = _RAND_158[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  mx2_5_4 = _RAND_159[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  mx2_5_5 = _RAND_160[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  mx2_5_6 = _RAND_161[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  mx2_5_7 = _RAND_162[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  mx2_6_0 = _RAND_163[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  mx2_6_1 = _RAND_164[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  mx2_6_2 = _RAND_165[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  mx2_6_3 = _RAND_166[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  mx2_6_4 = _RAND_167[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  mx2_6_5 = _RAND_168[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  mx2_6_6 = _RAND_169[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  mx2_6_7 = _RAND_170[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  mx2_7_0 = _RAND_171[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  mx2_7_1 = _RAND_172[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  mx2_7_2 = _RAND_173[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  mx2_7_3 = _RAND_174[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  mx2_7_4 = _RAND_175[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  mx2_7_5 = _RAND_176[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  mx2_7_6 = _RAND_177[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  mx2_7_7 = _RAND_178[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  ab2_0_0 = _RAND_179[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  ab2_0_1 = _RAND_180[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  ab2_0_2 = _RAND_181[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  ab2_0_3 = _RAND_182[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  ab2_0_4 = _RAND_183[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  ab2_0_5 = _RAND_184[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  ab2_0_6 = _RAND_185[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  ab2_0_7 = _RAND_186[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  ab2_1_0 = _RAND_187[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  ab2_1_1 = _RAND_188[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  ab2_1_2 = _RAND_189[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  ab2_1_3 = _RAND_190[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  ab2_1_4 = _RAND_191[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  ab2_1_5 = _RAND_192[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  ab2_1_6 = _RAND_193[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  ab2_1_7 = _RAND_194[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  ab2_2_0 = _RAND_195[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  ab2_2_1 = _RAND_196[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  ab2_2_2 = _RAND_197[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  ab2_2_3 = _RAND_198[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  ab2_2_4 = _RAND_199[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  ab2_2_5 = _RAND_200[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{`RANDOM}};
  ab2_2_6 = _RAND_201[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{`RANDOM}};
  ab2_2_7 = _RAND_202[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{`RANDOM}};
  ab2_3_0 = _RAND_203[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{`RANDOM}};
  ab2_3_1 = _RAND_204[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{`RANDOM}};
  ab2_3_2 = _RAND_205[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{`RANDOM}};
  ab2_3_3 = _RAND_206[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{`RANDOM}};
  ab2_3_4 = _RAND_207[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{`RANDOM}};
  ab2_3_5 = _RAND_208[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{`RANDOM}};
  ab2_3_6 = _RAND_209[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{`RANDOM}};
  ab2_3_7 = _RAND_210[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{`RANDOM}};
  ab2_4_0 = _RAND_211[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{`RANDOM}};
  ab2_4_1 = _RAND_212[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{`RANDOM}};
  ab2_4_2 = _RAND_213[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{`RANDOM}};
  ab2_4_3 = _RAND_214[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{`RANDOM}};
  ab2_4_4 = _RAND_215[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{`RANDOM}};
  ab2_4_5 = _RAND_216[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{`RANDOM}};
  ab2_4_6 = _RAND_217[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{`RANDOM}};
  ab2_4_7 = _RAND_218[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{`RANDOM}};
  ab2_5_0 = _RAND_219[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{`RANDOM}};
  ab2_5_1 = _RAND_220[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{`RANDOM}};
  ab2_5_2 = _RAND_221[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{`RANDOM}};
  ab2_5_3 = _RAND_222[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{`RANDOM}};
  ab2_5_4 = _RAND_223[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{`RANDOM}};
  ab2_5_5 = _RAND_224[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{`RANDOM}};
  ab2_5_6 = _RAND_225[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{`RANDOM}};
  ab2_5_7 = _RAND_226[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{`RANDOM}};
  ab2_6_0 = _RAND_227[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{`RANDOM}};
  ab2_6_1 = _RAND_228[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{`RANDOM}};
  ab2_6_2 = _RAND_229[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{`RANDOM}};
  ab2_6_3 = _RAND_230[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{`RANDOM}};
  ab2_6_4 = _RAND_231[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{`RANDOM}};
  ab2_6_5 = _RAND_232[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{`RANDOM}};
  ab2_6_6 = _RAND_233[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{`RANDOM}};
  ab2_6_7 = _RAND_234[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{`RANDOM}};
  ab2_7_0 = _RAND_235[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{`RANDOM}};
  ab2_7_1 = _RAND_236[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{`RANDOM}};
  ab2_7_2 = _RAND_237[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{`RANDOM}};
  ab2_7_3 = _RAND_238[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{`RANDOM}};
  ab2_7_4 = _RAND_239[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{`RANDOM}};
  ab2_7_5 = _RAND_240[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{`RANDOM}};
  ab2_7_6 = _RAND_241[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{`RANDOM}};
  ab2_7_7 = _RAND_242[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{`RANDOM}};
  tm8_0_0 = _RAND_243[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{`RANDOM}};
  tm8_0_1 = _RAND_244[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{`RANDOM}};
  tm8_0_2 = _RAND_245[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{`RANDOM}};
  tm8_0_3 = _RAND_246[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{`RANDOM}};
  tm8_0_4 = _RAND_247[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{`RANDOM}};
  tm8_0_5 = _RAND_248[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{`RANDOM}};
  tm8_0_6 = _RAND_249[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{`RANDOM}};
  tm8_0_7 = _RAND_250[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{`RANDOM}};
  tm8_1_0 = _RAND_251[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{`RANDOM}};
  tm8_1_1 = _RAND_252[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{`RANDOM}};
  tm8_1_2 = _RAND_253[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{`RANDOM}};
  tm8_1_3 = _RAND_254[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{`RANDOM}};
  tm8_1_4 = _RAND_255[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_256 = {1{`RANDOM}};
  tm8_1_5 = _RAND_256[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_257 = {1{`RANDOM}};
  tm8_1_6 = _RAND_257[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_258 = {1{`RANDOM}};
  tm8_1_7 = _RAND_258[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_259 = {1{`RANDOM}};
  tm8_2_0 = _RAND_259[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_260 = {1{`RANDOM}};
  tm8_2_1 = _RAND_260[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_261 = {1{`RANDOM}};
  tm8_2_2 = _RAND_261[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_262 = {1{`RANDOM}};
  tm8_2_3 = _RAND_262[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_263 = {1{`RANDOM}};
  tm8_2_4 = _RAND_263[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_264 = {1{`RANDOM}};
  tm8_2_5 = _RAND_264[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_265 = {1{`RANDOM}};
  tm8_2_6 = _RAND_265[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_266 = {1{`RANDOM}};
  tm8_2_7 = _RAND_266[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_267 = {1{`RANDOM}};
  tm8_3_0 = _RAND_267[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_268 = {1{`RANDOM}};
  tm8_3_1 = _RAND_268[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_269 = {1{`RANDOM}};
  tm8_3_2 = _RAND_269[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_270 = {1{`RANDOM}};
  tm8_3_3 = _RAND_270[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_271 = {1{`RANDOM}};
  tm8_3_4 = _RAND_271[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_272 = {1{`RANDOM}};
  tm8_3_5 = _RAND_272[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_273 = {1{`RANDOM}};
  tm8_3_6 = _RAND_273[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_274 = {1{`RANDOM}};
  tm8_3_7 = _RAND_274[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_275 = {1{`RANDOM}};
  tm9_0_0 = _RAND_275[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_276 = {1{`RANDOM}};
  tm9_0_1 = _RAND_276[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_277 = {1{`RANDOM}};
  tm9_0_2 = _RAND_277[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_278 = {1{`RANDOM}};
  tm9_0_3 = _RAND_278[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_279 = {1{`RANDOM}};
  tm9_0_4 = _RAND_279[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_280 = {1{`RANDOM}};
  tm9_0_5 = _RAND_280[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_281 = {1{`RANDOM}};
  tm9_0_6 = _RAND_281[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_282 = {1{`RANDOM}};
  tm9_0_7 = _RAND_282[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_283 = {1{`RANDOM}};
  tm9_1_0 = _RAND_283[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_284 = {1{`RANDOM}};
  tm9_1_1 = _RAND_284[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_285 = {1{`RANDOM}};
  tm9_1_2 = _RAND_285[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_286 = {1{`RANDOM}};
  tm9_1_3 = _RAND_286[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_287 = {1{`RANDOM}};
  tm9_1_4 = _RAND_287[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_288 = {1{`RANDOM}};
  tm9_1_5 = _RAND_288[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_289 = {1{`RANDOM}};
  tm9_1_6 = _RAND_289[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_290 = {1{`RANDOM}};
  tm9_1_7 = _RAND_290[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_291 = {1{`RANDOM}};
  tma_0_0 = _RAND_291[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_292 = {1{`RANDOM}};
  tma_0_1 = _RAND_292[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_293 = {1{`RANDOM}};
  tma_0_2 = _RAND_293[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_294 = {1{`RANDOM}};
  tma_0_3 = _RAND_294[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_295 = {1{`RANDOM}};
  tma_0_4 = _RAND_295[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_296 = {1{`RANDOM}};
  tma_0_5 = _RAND_296[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_297 = {1{`RANDOM}};
  tma_0_6 = _RAND_297[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_298 = {1{`RANDOM}};
  tma_0_7 = _RAND_298[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_299 = {1{`RANDOM}};
  tmb_0_0 = _RAND_299[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_300 = {1{`RANDOM}};
  tmb_0_1 = _RAND_300[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_301 = {1{`RANDOM}};
  tmb_0_2 = _RAND_301[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_302 = {1{`RANDOM}};
  tmb_0_3 = _RAND_302[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_303 = {1{`RANDOM}};
  tmb_0_4 = _RAND_303[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_304 = {1{`RANDOM}};
  tmb_0_5 = _RAND_304[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_305 = {1{`RANDOM}};
  tmb_0_6 = _RAND_305[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_306 = {1{`RANDOM}};
  tmb_0_7 = _RAND_306[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_307 = {1{`RANDOM}};
  tmc_0_0 = _RAND_307[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_308 = {1{`RANDOM}};
  tmc_0_1 = _RAND_308[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_309 = {1{`RANDOM}};
  tmc_0_2 = _RAND_309[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_310 = {1{`RANDOM}};
  tmc_0_3 = _RAND_310[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_311 = {1{`RANDOM}};
  tmc_0_4 = _RAND_311[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_312 = {1{`RANDOM}};
  tmc_0_5 = _RAND_312[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_313 = {1{`RANDOM}};
  tmc_0_6 = _RAND_313[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_314 = {1{`RANDOM}};
  tmc_0_7 = _RAND_314[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_315 = {1{`RANDOM}};
  best_0 = _RAND_315[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_316 = {1{`RANDOM}};
  best_1 = _RAND_316[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_317 = {1{`RANDOM}};
  best_2 = _RAND_317[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_318 = {1{`RANDOM}};
  best_3 = _RAND_318[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_319 = {1{`RANDOM}};
  best_4 = _RAND_319[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_320 = {1{`RANDOM}};
  best_5 = _RAND_320[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_321 = {1{`RANDOM}};
  best_6 = _RAND_321[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_322 = {1{`RANDOM}};
  best_7 = _RAND_322[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_323 = {1{`RANDOM}};
  bestBufe_0 = _RAND_323[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_324 = {1{`RANDOM}};
  bestBufe_1 = _RAND_324[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_325 = {1{`RANDOM}};
  bestBufe_2 = _RAND_325[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_326 = {1{`RANDOM}};
  bestBufe_3 = _RAND_326[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_327 = {1{`RANDOM}};
  bestBufe_4 = _RAND_327[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_328 = {1{`RANDOM}};
  bestBufe_5 = _RAND_328[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_329 = {1{`RANDOM}};
  bestBufe_6 = _RAND_329[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_330 = {1{`RANDOM}};
  bestBufe_7 = _RAND_330[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_331 = {1{`RANDOM}};
  r = _RAND_331[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_332 = {1{`RANDOM}};
  c = _RAND_332[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_333 = {1{`RANDOM}};
  BFbuf_e = _RAND_333[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_334 = {1{`RANDOM}};
  BFbuf_a = _RAND_334[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_335 = {1{`RANDOM}};
  load_i = _RAND_335[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_336 = {1{`RANDOM}};
  load_j = _RAND_336[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_337 = {1{`RANDOM}};
  doneLoading = _RAND_337[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_338 = {1{`RANDOM}};
  lastLoad = _RAND_338[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_339 = {1{`RANDOM}};
  prev_lo_i = _RAND_339[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_340 = {1{`RANDOM}};
  prev_lo_j = _RAND_340[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_341 = {1{`RANDOM}};
  prev_idx = _RAND_341[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_342 = {1{`RANDOM}};
  slcBuf_e = _RAND_342[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_343 = {1{`RANDOM}};
  slcBuf_a = _RAND_343[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_344 = {1{`RANDOM}};
  slcValid = _RAND_344[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_345 = {1{`RANDOM}};
  AEbuf_0_0_e = _RAND_345[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_346 = {1{`RANDOM}};
  AEbuf_0_0_a = _RAND_346[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_347 = {1{`RANDOM}};
  AEbuf_0_1_e = _RAND_347[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_348 = {1{`RANDOM}};
  AEbuf_0_1_a = _RAND_348[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_349 = {1{`RANDOM}};
  AEbuf_0_2_e = _RAND_349[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_350 = {1{`RANDOM}};
  AEbuf_0_2_a = _RAND_350[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_351 = {1{`RANDOM}};
  AEbuf_0_3_e = _RAND_351[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_352 = {1{`RANDOM}};
  AEbuf_0_3_a = _RAND_352[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_353 = {1{`RANDOM}};
  AEbuf_0_4_e = _RAND_353[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_354 = {1{`RANDOM}};
  AEbuf_0_4_a = _RAND_354[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_355 = {1{`RANDOM}};
  AEbuf_0_5_e = _RAND_355[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_356 = {1{`RANDOM}};
  AEbuf_0_5_a = _RAND_356[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_357 = {1{`RANDOM}};
  AEbuf_0_6_e = _RAND_357[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_358 = {1{`RANDOM}};
  AEbuf_0_6_a = _RAND_358[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_359 = {1{`RANDOM}};
  AEbuf_0_7_e = _RAND_359[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_360 = {1{`RANDOM}};
  AEbuf_0_7_a = _RAND_360[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_361 = {1{`RANDOM}};
  AEbuf_1_0_e = _RAND_361[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_362 = {1{`RANDOM}};
  AEbuf_1_0_a = _RAND_362[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_363 = {1{`RANDOM}};
  AEbuf_1_1_e = _RAND_363[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_364 = {1{`RANDOM}};
  AEbuf_1_1_a = _RAND_364[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_365 = {1{`RANDOM}};
  AEbuf_1_2_e = _RAND_365[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_366 = {1{`RANDOM}};
  AEbuf_1_2_a = _RAND_366[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_367 = {1{`RANDOM}};
  AEbuf_1_3_e = _RAND_367[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_368 = {1{`RANDOM}};
  AEbuf_1_3_a = _RAND_368[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_369 = {1{`RANDOM}};
  AEbuf_1_4_e = _RAND_369[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_370 = {1{`RANDOM}};
  AEbuf_1_4_a = _RAND_370[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_371 = {1{`RANDOM}};
  AEbuf_1_5_e = _RAND_371[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_372 = {1{`RANDOM}};
  AEbuf_1_5_a = _RAND_372[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_373 = {1{`RANDOM}};
  AEbuf_1_6_e = _RAND_373[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_374 = {1{`RANDOM}};
  AEbuf_1_6_a = _RAND_374[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_375 = {1{`RANDOM}};
  AEbuf_1_7_e = _RAND_375[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_376 = {1{`RANDOM}};
  AEbuf_1_7_a = _RAND_376[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_377 = {1{`RANDOM}};
  AEbuf_2_0_e = _RAND_377[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_378 = {1{`RANDOM}};
  AEbuf_2_0_a = _RAND_378[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_379 = {1{`RANDOM}};
  AEbuf_2_1_e = _RAND_379[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_380 = {1{`RANDOM}};
  AEbuf_2_1_a = _RAND_380[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_381 = {1{`RANDOM}};
  AEbuf_2_2_e = _RAND_381[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_382 = {1{`RANDOM}};
  AEbuf_2_2_a = _RAND_382[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_383 = {1{`RANDOM}};
  AEbuf_2_3_e = _RAND_383[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_384 = {1{`RANDOM}};
  AEbuf_2_3_a = _RAND_384[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_385 = {1{`RANDOM}};
  AEbuf_2_4_e = _RAND_385[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_386 = {1{`RANDOM}};
  AEbuf_2_4_a = _RAND_386[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_387 = {1{`RANDOM}};
  AEbuf_2_5_e = _RAND_387[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_388 = {1{`RANDOM}};
  AEbuf_2_5_a = _RAND_388[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_389 = {1{`RANDOM}};
  AEbuf_2_6_e = _RAND_389[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_390 = {1{`RANDOM}};
  AEbuf_2_6_a = _RAND_390[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_391 = {1{`RANDOM}};
  AEbuf_2_7_e = _RAND_391[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_392 = {1{`RANDOM}};
  AEbuf_2_7_a = _RAND_392[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_393 = {1{`RANDOM}};
  AEbuf_3_0_e = _RAND_393[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_394 = {1{`RANDOM}};
  AEbuf_3_0_a = _RAND_394[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_395 = {1{`RANDOM}};
  AEbuf_3_1_e = _RAND_395[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_396 = {1{`RANDOM}};
  AEbuf_3_1_a = _RAND_396[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_397 = {1{`RANDOM}};
  AEbuf_3_2_e = _RAND_397[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_398 = {1{`RANDOM}};
  AEbuf_3_2_a = _RAND_398[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_399 = {1{`RANDOM}};
  AEbuf_3_3_e = _RAND_399[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_400 = {1{`RANDOM}};
  AEbuf_3_3_a = _RAND_400[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_401 = {1{`RANDOM}};
  AEbuf_3_4_e = _RAND_401[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_402 = {1{`RANDOM}};
  AEbuf_3_4_a = _RAND_402[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_403 = {1{`RANDOM}};
  AEbuf_3_5_e = _RAND_403[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_404 = {1{`RANDOM}};
  AEbuf_3_5_a = _RAND_404[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_405 = {1{`RANDOM}};
  AEbuf_3_6_e = _RAND_405[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_406 = {1{`RANDOM}};
  AEbuf_3_6_a = _RAND_406[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_407 = {1{`RANDOM}};
  AEbuf_3_7_e = _RAND_407[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_408 = {1{`RANDOM}};
  AEbuf_3_7_a = _RAND_408[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_409 = {1{`RANDOM}};
  AEbuf_4_0_e = _RAND_409[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_410 = {1{`RANDOM}};
  AEbuf_4_0_a = _RAND_410[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_411 = {1{`RANDOM}};
  AEbuf_4_1_e = _RAND_411[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_412 = {1{`RANDOM}};
  AEbuf_4_1_a = _RAND_412[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_413 = {1{`RANDOM}};
  AEbuf_4_2_e = _RAND_413[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_414 = {1{`RANDOM}};
  AEbuf_4_2_a = _RAND_414[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_415 = {1{`RANDOM}};
  AEbuf_4_3_e = _RAND_415[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_416 = {1{`RANDOM}};
  AEbuf_4_3_a = _RAND_416[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_417 = {1{`RANDOM}};
  AEbuf_4_4_e = _RAND_417[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_418 = {1{`RANDOM}};
  AEbuf_4_4_a = _RAND_418[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_419 = {1{`RANDOM}};
  AEbuf_4_5_e = _RAND_419[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_420 = {1{`RANDOM}};
  AEbuf_4_5_a = _RAND_420[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_421 = {1{`RANDOM}};
  AEbuf_4_6_e = _RAND_421[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_422 = {1{`RANDOM}};
  AEbuf_4_6_a = _RAND_422[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_423 = {1{`RANDOM}};
  AEbuf_4_7_e = _RAND_423[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_424 = {1{`RANDOM}};
  AEbuf_4_7_a = _RAND_424[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_425 = {1{`RANDOM}};
  AEbuf_5_0_e = _RAND_425[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_426 = {1{`RANDOM}};
  AEbuf_5_0_a = _RAND_426[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_427 = {1{`RANDOM}};
  AEbuf_5_1_e = _RAND_427[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_428 = {1{`RANDOM}};
  AEbuf_5_1_a = _RAND_428[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_429 = {1{`RANDOM}};
  AEbuf_5_2_e = _RAND_429[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_430 = {1{`RANDOM}};
  AEbuf_5_2_a = _RAND_430[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_431 = {1{`RANDOM}};
  AEbuf_5_3_e = _RAND_431[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_432 = {1{`RANDOM}};
  AEbuf_5_3_a = _RAND_432[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_433 = {1{`RANDOM}};
  AEbuf_5_4_e = _RAND_433[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_434 = {1{`RANDOM}};
  AEbuf_5_4_a = _RAND_434[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_435 = {1{`RANDOM}};
  AEbuf_5_5_e = _RAND_435[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_436 = {1{`RANDOM}};
  AEbuf_5_5_a = _RAND_436[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_437 = {1{`RANDOM}};
  AEbuf_5_6_e = _RAND_437[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_438 = {1{`RANDOM}};
  AEbuf_5_6_a = _RAND_438[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_439 = {1{`RANDOM}};
  AEbuf_5_7_e = _RAND_439[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_440 = {1{`RANDOM}};
  AEbuf_5_7_a = _RAND_440[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_441 = {1{`RANDOM}};
  AEbuf_6_0_e = _RAND_441[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_442 = {1{`RANDOM}};
  AEbuf_6_0_a = _RAND_442[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_443 = {1{`RANDOM}};
  AEbuf_6_1_e = _RAND_443[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_444 = {1{`RANDOM}};
  AEbuf_6_1_a = _RAND_444[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_445 = {1{`RANDOM}};
  AEbuf_6_2_e = _RAND_445[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_446 = {1{`RANDOM}};
  AEbuf_6_2_a = _RAND_446[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_447 = {1{`RANDOM}};
  AEbuf_6_3_e = _RAND_447[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_448 = {1{`RANDOM}};
  AEbuf_6_3_a = _RAND_448[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_449 = {1{`RANDOM}};
  AEbuf_6_4_e = _RAND_449[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_450 = {1{`RANDOM}};
  AEbuf_6_4_a = _RAND_450[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_451 = {1{`RANDOM}};
  AEbuf_6_5_e = _RAND_451[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_452 = {1{`RANDOM}};
  AEbuf_6_5_a = _RAND_452[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_453 = {1{`RANDOM}};
  AEbuf_6_6_e = _RAND_453[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_454 = {1{`RANDOM}};
  AEbuf_6_6_a = _RAND_454[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_455 = {1{`RANDOM}};
  AEbuf_6_7_e = _RAND_455[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_456 = {1{`RANDOM}};
  AEbuf_6_7_a = _RAND_456[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_457 = {1{`RANDOM}};
  AEbuf_7_0_e = _RAND_457[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_458 = {1{`RANDOM}};
  AEbuf_7_0_a = _RAND_458[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_459 = {1{`RANDOM}};
  AEbuf_7_1_e = _RAND_459[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_460 = {1{`RANDOM}};
  AEbuf_7_1_a = _RAND_460[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_461 = {1{`RANDOM}};
  AEbuf_7_2_e = _RAND_461[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_462 = {1{`RANDOM}};
  AEbuf_7_2_a = _RAND_462[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_463 = {1{`RANDOM}};
  AEbuf_7_3_e = _RAND_463[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_464 = {1{`RANDOM}};
  AEbuf_7_3_a = _RAND_464[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_465 = {1{`RANDOM}};
  AEbuf_7_4_e = _RAND_465[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_466 = {1{`RANDOM}};
  AEbuf_7_4_a = _RAND_466[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_467 = {1{`RANDOM}};
  AEbuf_7_5_e = _RAND_467[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_468 = {1{`RANDOM}};
  AEbuf_7_5_a = _RAND_468[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_469 = {1{`RANDOM}};
  AEbuf_7_6_e = _RAND_469[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_470 = {1{`RANDOM}};
  AEbuf_7_6_a = _RAND_470[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_471 = {1{`RANDOM}};
  AEbuf_7_7_e = _RAND_471[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_472 = {1{`RANDOM}};
  AEbuf_7_7_a = _RAND_472[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_473 = {1{`RANDOM}};
  _T_405 = _RAND_473[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_474 = {1{`RANDOM}};
  _T_406 = _RAND_474[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_475 = {1{`RANDOM}};
  _T_407 = _RAND_475[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_476 = {1{`RANDOM}};
  _T_408 = _RAND_476[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_477 = {1{`RANDOM}};
  _T_409 = _RAND_477[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_478 = {1{`RANDOM}};
  _T_410 = _RAND_478[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_479 = {1{`RANDOM}};
  _T_411 = _RAND_479[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_480 = {1{`RANDOM}};
  _T_412 = _RAND_480[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_481 = {1{`RANDOM}};
  _T_413 = _RAND_481[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_482 = {1{`RANDOM}};
  _T_414 = _RAND_482[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_483 = {1{`RANDOM}};
  _T_415 = _RAND_483[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_484 = {1{`RANDOM}};
  _T_416 = _RAND_484[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_485 = {1{`RANDOM}};
  _T_417 = _RAND_485[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_486 = {1{`RANDOM}};
  _T_418 = _RAND_486[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_487 = {1{`RANDOM}};
  _T_421 = _RAND_487[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_488 = {1{`RANDOM}};
  _T_422 = _RAND_488[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_489 = {1{`RANDOM}};
  _T_423 = _RAND_489[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_490 = {1{`RANDOM}};
  _T_424 = _RAND_490[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_491 = {1{`RANDOM}};
  _T_425 = _RAND_491[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_492 = {1{`RANDOM}};
  _T_426 = _RAND_492[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_493 = {1{`RANDOM}};
  _T_427 = _RAND_493[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_494 = {1{`RANDOM}};
  _T_428 = _RAND_494[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_495 = {1{`RANDOM}};
  _T_429 = _RAND_495[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_496 = {1{`RANDOM}};
  _T_430 = _RAND_496[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_497 = {1{`RANDOM}};
  _T_431 = _RAND_497[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_498 = {1{`RANDOM}};
  _T_432 = _RAND_498[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_499 = {1{`RANDOM}};
  _T_433 = _RAND_499[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_500 = {1{`RANDOM}};
  _T_434 = _RAND_500[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_501 = {1{`RANDOM}};
  _T_437 = _RAND_501[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_502 = {1{`RANDOM}};
  _T_438 = _RAND_502[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_503 = {1{`RANDOM}};
  _T_439 = _RAND_503[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_504 = {1{`RANDOM}};
  _T_440 = _RAND_504[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_505 = {1{`RANDOM}};
  _T_441 = _RAND_505[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_506 = {1{`RANDOM}};
  _T_442 = _RAND_506[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_507 = {1{`RANDOM}};
  _T_443 = _RAND_507[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_508 = {1{`RANDOM}};
  _T_444 = _RAND_508[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_509 = {1{`RANDOM}};
  _T_445 = _RAND_509[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_510 = {1{`RANDOM}};
  _T_446 = _RAND_510[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_511 = {1{`RANDOM}};
  _T_447 = _RAND_511[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_512 = {1{`RANDOM}};
  _T_448 = _RAND_512[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(AE_0_0__T_9_en & AE_0_0__T_9_mask) begin
      AE_0_0[AE_0_0__T_9_addr] <= AE_0_0__T_9_data; // @[loaf.scala 147:67]
    end
    if(AE_0_1__T_15_en & AE_0_1__T_15_mask) begin
      AE_0_1[AE_0_1__T_15_addr] <= AE_0_1__T_15_data; // @[loaf.scala 147:67]
    end
    if(AE_0_2__T_21_en & AE_0_2__T_21_mask) begin
      AE_0_2[AE_0_2__T_21_addr] <= AE_0_2__T_21_data; // @[loaf.scala 147:67]
    end
    if(AE_0_3__T_27_en & AE_0_3__T_27_mask) begin
      AE_0_3[AE_0_3__T_27_addr] <= AE_0_3__T_27_data; // @[loaf.scala 147:67]
    end
    if(AE_0_4__T_33_en & AE_0_4__T_33_mask) begin
      AE_0_4[AE_0_4__T_33_addr] <= AE_0_4__T_33_data; // @[loaf.scala 147:67]
    end
    if(AE_0_5__T_39_en & AE_0_5__T_39_mask) begin
      AE_0_5[AE_0_5__T_39_addr] <= AE_0_5__T_39_data; // @[loaf.scala 147:67]
    end
    if(AE_0_6__T_45_en & AE_0_6__T_45_mask) begin
      AE_0_6[AE_0_6__T_45_addr] <= AE_0_6__T_45_data; // @[loaf.scala 147:67]
    end
    if(AE_0_7__T_51_en & AE_0_7__T_51_mask) begin
      AE_0_7[AE_0_7__T_51_addr] <= AE_0_7__T_51_data; // @[loaf.scala 147:67]
    end
    if(AE_1_0__T_57_en & AE_1_0__T_57_mask) begin
      AE_1_0[AE_1_0__T_57_addr] <= AE_1_0__T_57_data; // @[loaf.scala 147:67]
    end
    if(AE_1_1__T_63_en & AE_1_1__T_63_mask) begin
      AE_1_1[AE_1_1__T_63_addr] <= AE_1_1__T_63_data; // @[loaf.scala 147:67]
    end
    if(AE_1_2__T_69_en & AE_1_2__T_69_mask) begin
      AE_1_2[AE_1_2__T_69_addr] <= AE_1_2__T_69_data; // @[loaf.scala 147:67]
    end
    if(AE_1_3__T_75_en & AE_1_3__T_75_mask) begin
      AE_1_3[AE_1_3__T_75_addr] <= AE_1_3__T_75_data; // @[loaf.scala 147:67]
    end
    if(AE_1_4__T_81_en & AE_1_4__T_81_mask) begin
      AE_1_4[AE_1_4__T_81_addr] <= AE_1_4__T_81_data; // @[loaf.scala 147:67]
    end
    if(AE_1_5__T_87_en & AE_1_5__T_87_mask) begin
      AE_1_5[AE_1_5__T_87_addr] <= AE_1_5__T_87_data; // @[loaf.scala 147:67]
    end
    if(AE_1_6__T_93_en & AE_1_6__T_93_mask) begin
      AE_1_6[AE_1_6__T_93_addr] <= AE_1_6__T_93_data; // @[loaf.scala 147:67]
    end
    if(AE_1_7__T_99_en & AE_1_7__T_99_mask) begin
      AE_1_7[AE_1_7__T_99_addr] <= AE_1_7__T_99_data; // @[loaf.scala 147:67]
    end
    if(AE_2_0__T_105_en & AE_2_0__T_105_mask) begin
      AE_2_0[AE_2_0__T_105_addr] <= AE_2_0__T_105_data; // @[loaf.scala 147:67]
    end
    if(AE_2_1__T_111_en & AE_2_1__T_111_mask) begin
      AE_2_1[AE_2_1__T_111_addr] <= AE_2_1__T_111_data; // @[loaf.scala 147:67]
    end
    if(AE_2_2__T_117_en & AE_2_2__T_117_mask) begin
      AE_2_2[AE_2_2__T_117_addr] <= AE_2_2__T_117_data; // @[loaf.scala 147:67]
    end
    if(AE_2_3__T_123_en & AE_2_3__T_123_mask) begin
      AE_2_3[AE_2_3__T_123_addr] <= AE_2_3__T_123_data; // @[loaf.scala 147:67]
    end
    if(AE_2_4__T_129_en & AE_2_4__T_129_mask) begin
      AE_2_4[AE_2_4__T_129_addr] <= AE_2_4__T_129_data; // @[loaf.scala 147:67]
    end
    if(AE_2_5__T_135_en & AE_2_5__T_135_mask) begin
      AE_2_5[AE_2_5__T_135_addr] <= AE_2_5__T_135_data; // @[loaf.scala 147:67]
    end
    if(AE_2_6__T_141_en & AE_2_6__T_141_mask) begin
      AE_2_6[AE_2_6__T_141_addr] <= AE_2_6__T_141_data; // @[loaf.scala 147:67]
    end
    if(AE_2_7__T_147_en & AE_2_7__T_147_mask) begin
      AE_2_7[AE_2_7__T_147_addr] <= AE_2_7__T_147_data; // @[loaf.scala 147:67]
    end
    if(AE_3_0__T_153_en & AE_3_0__T_153_mask) begin
      AE_3_0[AE_3_0__T_153_addr] <= AE_3_0__T_153_data; // @[loaf.scala 147:67]
    end
    if(AE_3_1__T_159_en & AE_3_1__T_159_mask) begin
      AE_3_1[AE_3_1__T_159_addr] <= AE_3_1__T_159_data; // @[loaf.scala 147:67]
    end
    if(AE_3_2__T_165_en & AE_3_2__T_165_mask) begin
      AE_3_2[AE_3_2__T_165_addr] <= AE_3_2__T_165_data; // @[loaf.scala 147:67]
    end
    if(AE_3_3__T_171_en & AE_3_3__T_171_mask) begin
      AE_3_3[AE_3_3__T_171_addr] <= AE_3_3__T_171_data; // @[loaf.scala 147:67]
    end
    if(AE_3_4__T_177_en & AE_3_4__T_177_mask) begin
      AE_3_4[AE_3_4__T_177_addr] <= AE_3_4__T_177_data; // @[loaf.scala 147:67]
    end
    if(AE_3_5__T_183_en & AE_3_5__T_183_mask) begin
      AE_3_5[AE_3_5__T_183_addr] <= AE_3_5__T_183_data; // @[loaf.scala 147:67]
    end
    if(AE_3_6__T_189_en & AE_3_6__T_189_mask) begin
      AE_3_6[AE_3_6__T_189_addr] <= AE_3_6__T_189_data; // @[loaf.scala 147:67]
    end
    if(AE_3_7__T_195_en & AE_3_7__T_195_mask) begin
      AE_3_7[AE_3_7__T_195_addr] <= AE_3_7__T_195_data; // @[loaf.scala 147:67]
    end
    if(AE_4_0__T_201_en & AE_4_0__T_201_mask) begin
      AE_4_0[AE_4_0__T_201_addr] <= AE_4_0__T_201_data; // @[loaf.scala 147:67]
    end
    if(AE_4_1__T_207_en & AE_4_1__T_207_mask) begin
      AE_4_1[AE_4_1__T_207_addr] <= AE_4_1__T_207_data; // @[loaf.scala 147:67]
    end
    if(AE_4_2__T_213_en & AE_4_2__T_213_mask) begin
      AE_4_2[AE_4_2__T_213_addr] <= AE_4_2__T_213_data; // @[loaf.scala 147:67]
    end
    if(AE_4_3__T_219_en & AE_4_3__T_219_mask) begin
      AE_4_3[AE_4_3__T_219_addr] <= AE_4_3__T_219_data; // @[loaf.scala 147:67]
    end
    if(AE_4_4__T_225_en & AE_4_4__T_225_mask) begin
      AE_4_4[AE_4_4__T_225_addr] <= AE_4_4__T_225_data; // @[loaf.scala 147:67]
    end
    if(AE_4_5__T_231_en & AE_4_5__T_231_mask) begin
      AE_4_5[AE_4_5__T_231_addr] <= AE_4_5__T_231_data; // @[loaf.scala 147:67]
    end
    if(AE_4_6__T_237_en & AE_4_6__T_237_mask) begin
      AE_4_6[AE_4_6__T_237_addr] <= AE_4_6__T_237_data; // @[loaf.scala 147:67]
    end
    if(AE_4_7__T_243_en & AE_4_7__T_243_mask) begin
      AE_4_7[AE_4_7__T_243_addr] <= AE_4_7__T_243_data; // @[loaf.scala 147:67]
    end
    if(AE_5_0__T_249_en & AE_5_0__T_249_mask) begin
      AE_5_0[AE_5_0__T_249_addr] <= AE_5_0__T_249_data; // @[loaf.scala 147:67]
    end
    if(AE_5_1__T_255_en & AE_5_1__T_255_mask) begin
      AE_5_1[AE_5_1__T_255_addr] <= AE_5_1__T_255_data; // @[loaf.scala 147:67]
    end
    if(AE_5_2__T_261_en & AE_5_2__T_261_mask) begin
      AE_5_2[AE_5_2__T_261_addr] <= AE_5_2__T_261_data; // @[loaf.scala 147:67]
    end
    if(AE_5_3__T_267_en & AE_5_3__T_267_mask) begin
      AE_5_3[AE_5_3__T_267_addr] <= AE_5_3__T_267_data; // @[loaf.scala 147:67]
    end
    if(AE_5_4__T_273_en & AE_5_4__T_273_mask) begin
      AE_5_4[AE_5_4__T_273_addr] <= AE_5_4__T_273_data; // @[loaf.scala 147:67]
    end
    if(AE_5_5__T_279_en & AE_5_5__T_279_mask) begin
      AE_5_5[AE_5_5__T_279_addr] <= AE_5_5__T_279_data; // @[loaf.scala 147:67]
    end
    if(AE_5_6__T_285_en & AE_5_6__T_285_mask) begin
      AE_5_6[AE_5_6__T_285_addr] <= AE_5_6__T_285_data; // @[loaf.scala 147:67]
    end
    if(AE_5_7__T_291_en & AE_5_7__T_291_mask) begin
      AE_5_7[AE_5_7__T_291_addr] <= AE_5_7__T_291_data; // @[loaf.scala 147:67]
    end
    if(AE_6_0__T_297_en & AE_6_0__T_297_mask) begin
      AE_6_0[AE_6_0__T_297_addr] <= AE_6_0__T_297_data; // @[loaf.scala 147:67]
    end
    if(AE_6_1__T_303_en & AE_6_1__T_303_mask) begin
      AE_6_1[AE_6_1__T_303_addr] <= AE_6_1__T_303_data; // @[loaf.scala 147:67]
    end
    if(AE_6_2__T_309_en & AE_6_2__T_309_mask) begin
      AE_6_2[AE_6_2__T_309_addr] <= AE_6_2__T_309_data; // @[loaf.scala 147:67]
    end
    if(AE_6_3__T_315_en & AE_6_3__T_315_mask) begin
      AE_6_3[AE_6_3__T_315_addr] <= AE_6_3__T_315_data; // @[loaf.scala 147:67]
    end
    if(AE_6_4__T_321_en & AE_6_4__T_321_mask) begin
      AE_6_4[AE_6_4__T_321_addr] <= AE_6_4__T_321_data; // @[loaf.scala 147:67]
    end
    if(AE_6_5__T_327_en & AE_6_5__T_327_mask) begin
      AE_6_5[AE_6_5__T_327_addr] <= AE_6_5__T_327_data; // @[loaf.scala 147:67]
    end
    if(AE_6_6__T_333_en & AE_6_6__T_333_mask) begin
      AE_6_6[AE_6_6__T_333_addr] <= AE_6_6__T_333_data; // @[loaf.scala 147:67]
    end
    if(AE_6_7__T_339_en & AE_6_7__T_339_mask) begin
      AE_6_7[AE_6_7__T_339_addr] <= AE_6_7__T_339_data; // @[loaf.scala 147:67]
    end
    if(AE_7_0__T_345_en & AE_7_0__T_345_mask) begin
      AE_7_0[AE_7_0__T_345_addr] <= AE_7_0__T_345_data; // @[loaf.scala 147:67]
    end
    if(AE_7_1__T_351_en & AE_7_1__T_351_mask) begin
      AE_7_1[AE_7_1__T_351_addr] <= AE_7_1__T_351_data; // @[loaf.scala 147:67]
    end
    if(AE_7_2__T_357_en & AE_7_2__T_357_mask) begin
      AE_7_2[AE_7_2__T_357_addr] <= AE_7_2__T_357_data; // @[loaf.scala 147:67]
    end
    if(AE_7_3__T_363_en & AE_7_3__T_363_mask) begin
      AE_7_3[AE_7_3__T_363_addr] <= AE_7_3__T_363_data; // @[loaf.scala 147:67]
    end
    if(AE_7_4__T_369_en & AE_7_4__T_369_mask) begin
      AE_7_4[AE_7_4__T_369_addr] <= AE_7_4__T_369_data; // @[loaf.scala 147:67]
    end
    if(AE_7_5__T_375_en & AE_7_5__T_375_mask) begin
      AE_7_5[AE_7_5__T_375_addr] <= AE_7_5__T_375_data; // @[loaf.scala 147:67]
    end
    if(AE_7_6__T_381_en & AE_7_6__T_381_mask) begin
      AE_7_6[AE_7_6__T_381_addr] <= AE_7_6__T_381_data; // @[loaf.scala 147:67]
    end
    if(AE_7_7__T_387_en & AE_7_7__T_387_mask) begin
      AE_7_7[AE_7_7__T_387_addr] <= AE_7_7__T_387_data; // @[loaf.scala 147:67]
    end
    if (reset) begin
      islice <= 9'h0;
    end else begin
      if (_T_451) begin
        if (_T_452) begin
          if (_T_463) begin
            if (_T_466) begin
              if (!(_T_2102)) begin
                if (!(_T_2105)) begin
                  if (_T_2108) begin
                    islice <= _T_2110;
                  end else begin
                    islice <= 9'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      done <= 1'h0;
    end else begin
      if (_T_451) begin
        if (_T_452) begin
          if (_T_463) begin
            if (phase) begin
              if (_T_2139) begin
                done <= 1'h1;
              end
            end
          end
        end else begin
          if (doneLoading) begin
            done <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      phase <= 1'h0;
    end else begin
      if (_T_451) begin
        if (_T_452) begin
          if (_T_463) begin
            if (_T_466) begin
              if (!(_T_2102)) begin
                if (!(_T_2105)) begin
                  if (!(_T_2108)) begin
                    phase <= 1'h1;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            if (_T_454) begin
              if (2'h0 == r) begin
                offCLs_0_0 <= io_off_bits_0;
              end
            end
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            if (_T_454) begin
              if (2'h0 == r) begin
                offCLs_0_1 <= io_off_bits_1;
              end
            end
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            if (_T_454) begin
              if (2'h0 == r) begin
                offCLs_0_2 <= io_off_bits_2;
              end
            end
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            if (_T_454) begin
              if (2'h0 == r) begin
                offCLs_0_3 <= io_off_bits_3;
              end
            end
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            if (_T_454) begin
              if (2'h0 == r) begin
                offCLs_0_4 <= io_off_bits_4;
              end
            end
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            if (_T_454) begin
              if (2'h0 == r) begin
                offCLs_0_5 <= io_off_bits_5;
              end
            end
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            if (_T_454) begin
              if (2'h0 == r) begin
                offCLs_0_6 <= io_off_bits_6;
              end
            end
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            if (_T_454) begin
              if (2'h0 == r) begin
                offCLs_0_7 <= io_off_bits_7;
              end
            end
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            if (_T_454) begin
              if (2'h1 == r) begin
                offCLs_1_0 <= io_off_bits_0;
              end
            end
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            if (_T_454) begin
              if (2'h1 == r) begin
                offCLs_1_1 <= io_off_bits_1;
              end
            end
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            if (_T_454) begin
              if (2'h1 == r) begin
                offCLs_1_2 <= io_off_bits_2;
              end
            end
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            if (_T_454) begin
              if (2'h1 == r) begin
                offCLs_1_3 <= io_off_bits_3;
              end
            end
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            if (_T_454) begin
              if (2'h1 == r) begin
                offCLs_1_4 <= io_off_bits_4;
              end
            end
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            if (_T_454) begin
              if (2'h1 == r) begin
                offCLs_1_5 <= io_off_bits_5;
              end
            end
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            if (_T_454) begin
              if (2'h1 == r) begin
                offCLs_1_6 <= io_off_bits_6;
              end
            end
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            if (_T_454) begin
              if (2'h1 == r) begin
                offCLs_1_7 <= io_off_bits_7;
              end
            end
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            if (_T_454) begin
              if (2'h2 == r) begin
                offCLs_2_0 <= io_off_bits_0;
              end
            end
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            if (_T_454) begin
              if (2'h2 == r) begin
                offCLs_2_1 <= io_off_bits_1;
              end
            end
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            if (_T_454) begin
              if (2'h2 == r) begin
                offCLs_2_2 <= io_off_bits_2;
              end
            end
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            if (_T_454) begin
              if (2'h2 == r) begin
                offCLs_2_3 <= io_off_bits_3;
              end
            end
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            if (_T_454) begin
              if (2'h2 == r) begin
                offCLs_2_4 <= io_off_bits_4;
              end
            end
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            if (_T_454) begin
              if (2'h2 == r) begin
                offCLs_2_5 <= io_off_bits_5;
              end
            end
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            if (_T_454) begin
              if (2'h2 == r) begin
                offCLs_2_6 <= io_off_bits_6;
              end
            end
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            if (_T_454) begin
              if (2'h2 == r) begin
                offCLs_2_7 <= io_off_bits_7;
              end
            end
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            if (_T_454) begin
              if (2'h3 == r) begin
                offCLs_3_0 <= io_off_bits_0;
              end
            end
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            if (_T_454) begin
              if (2'h3 == r) begin
                offCLs_3_1 <= io_off_bits_1;
              end
            end
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            if (_T_454) begin
              if (2'h3 == r) begin
                offCLs_3_2 <= io_off_bits_2;
              end
            end
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            if (_T_454) begin
              if (2'h3 == r) begin
                offCLs_3_3 <= io_off_bits_3;
              end
            end
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            if (_T_454) begin
              if (2'h3 == r) begin
                offCLs_3_4 <= io_off_bits_4;
              end
            end
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            if (_T_454) begin
              if (2'h3 == r) begin
                offCLs_3_5 <= io_off_bits_5;
              end
            end
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            if (_T_454) begin
              if (2'h3 == r) begin
                offCLs_3_6 <= io_off_bits_6;
              end
            end
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            if (_T_454) begin
              if (2'h3 == r) begin
                offCLs_3_7 <= io_off_bits_7;
              end
            end
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            if (_T_454) begin
              o1_0 <= io_off_bits_0;
            end else begin
              if (2'h3 == r) begin
                o1_0 <= offCLs_3_0;
              end else begin
                if (2'h2 == r) begin
                  o1_0 <= offCLs_2_0;
                end else begin
                  if (2'h1 == r) begin
                    o1_0 <= offCLs_1_0;
                  end else begin
                    o1_0 <= offCLs_0_0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            if (_T_454) begin
              o1_1 <= io_off_bits_1;
            end else begin
              if (2'h3 == r) begin
                o1_1 <= offCLs_3_1;
              end else begin
                if (2'h2 == r) begin
                  o1_1 <= offCLs_2_1;
                end else begin
                  if (2'h1 == r) begin
                    o1_1 <= offCLs_1_1;
                  end else begin
                    o1_1 <= offCLs_0_1;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            if (_T_454) begin
              o1_2 <= io_off_bits_2;
            end else begin
              if (2'h3 == r) begin
                o1_2 <= offCLs_3_2;
              end else begin
                if (2'h2 == r) begin
                  o1_2 <= offCLs_2_2;
                end else begin
                  if (2'h1 == r) begin
                    o1_2 <= offCLs_1_2;
                  end else begin
                    o1_2 <= offCLs_0_2;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            if (_T_454) begin
              o1_3 <= io_off_bits_3;
            end else begin
              if (2'h3 == r) begin
                o1_3 <= offCLs_3_3;
              end else begin
                if (2'h2 == r) begin
                  o1_3 <= offCLs_2_3;
                end else begin
                  if (2'h1 == r) begin
                    o1_3 <= offCLs_1_3;
                  end else begin
                    o1_3 <= offCLs_0_3;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            if (_T_454) begin
              o1_4 <= io_off_bits_4;
            end else begin
              if (2'h3 == r) begin
                o1_4 <= offCLs_3_4;
              end else begin
                if (2'h2 == r) begin
                  o1_4 <= offCLs_2_4;
                end else begin
                  if (2'h1 == r) begin
                    o1_4 <= offCLs_1_4;
                  end else begin
                    o1_4 <= offCLs_0_4;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            if (_T_454) begin
              o1_5 <= io_off_bits_5;
            end else begin
              if (2'h3 == r) begin
                o1_5 <= offCLs_3_5;
              end else begin
                if (2'h2 == r) begin
                  o1_5 <= offCLs_2_5;
                end else begin
                  if (2'h1 == r) begin
                    o1_5 <= offCLs_1_5;
                  end else begin
                    o1_5 <= offCLs_0_5;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            if (_T_454) begin
              o1_6 <= io_off_bits_6;
            end else begin
              if (2'h3 == r) begin
                o1_6 <= offCLs_3_6;
              end else begin
                if (2'h2 == r) begin
                  o1_6 <= offCLs_2_6;
                end else begin
                  if (2'h1 == r) begin
                    o1_6 <= offCLs_1_6;
                  end else begin
                    o1_6 <= offCLs_0_6;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            if (_T_454) begin
              o1_7 <= io_off_bits_7;
            end else begin
              if (2'h3 == r) begin
                o1_7 <= offCLs_3_7;
              end else begin
                if (2'h2 == r) begin
                  o1_7 <= offCLs_2_7;
                end else begin
                  if (2'h1 == r) begin
                    o1_7 <= offCLs_1_7;
                  end else begin
                    o1_7 <= offCLs_0_7;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          o2_0 <= o1_0;
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          o2_1 <= o1_1;
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          o2_2 <= o1_2;
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          o2_3 <= o1_3;
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          o2_4 <= o1_4;
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          o2_5 <= o1_5;
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          o2_6 <= o1_6;
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          o2_7 <= o1_7;
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1196) begin
            mx2_0_0 <= BFbuf_e;
          end else begin
            mx2_0_0 <= AEbuf_0_0_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1309) begin
            mx2_0_1 <= BFbuf_e;
          end else begin
            mx2_0_1 <= AEbuf_0_1_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1422) begin
            mx2_0_2 <= BFbuf_e;
          end else begin
            mx2_0_2 <= AEbuf_0_2_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1535) begin
            mx2_0_3 <= BFbuf_e;
          end else begin
            mx2_0_3 <= AEbuf_0_3_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1648) begin
            mx2_0_4 <= BFbuf_e;
          end else begin
            mx2_0_4 <= AEbuf_0_4_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1761) begin
            mx2_0_5 <= BFbuf_e;
          end else begin
            mx2_0_5 <= AEbuf_0_5_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1874) begin
            mx2_0_6 <= BFbuf_e;
          end else begin
            mx2_0_6 <= AEbuf_0_6_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1987) begin
            mx2_0_7 <= BFbuf_e;
          end else begin
            mx2_0_7 <= AEbuf_0_7_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1208) begin
            mx2_1_0 <= BFbuf_e;
          end else begin
            mx2_1_0 <= AEbuf_1_0_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1321) begin
            mx2_1_1 <= BFbuf_e;
          end else begin
            mx2_1_1 <= AEbuf_1_1_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1434) begin
            mx2_1_2 <= BFbuf_e;
          end else begin
            mx2_1_2 <= AEbuf_1_2_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1547) begin
            mx2_1_3 <= BFbuf_e;
          end else begin
            mx2_1_3 <= AEbuf_1_3_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1660) begin
            mx2_1_4 <= BFbuf_e;
          end else begin
            mx2_1_4 <= AEbuf_1_4_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1773) begin
            mx2_1_5 <= BFbuf_e;
          end else begin
            mx2_1_5 <= AEbuf_1_5_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1886) begin
            mx2_1_6 <= BFbuf_e;
          end else begin
            mx2_1_6 <= AEbuf_1_6_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1999) begin
            mx2_1_7 <= BFbuf_e;
          end else begin
            mx2_1_7 <= AEbuf_1_7_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1220) begin
            mx2_2_0 <= BFbuf_e;
          end else begin
            mx2_2_0 <= AEbuf_2_0_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1333) begin
            mx2_2_1 <= BFbuf_e;
          end else begin
            mx2_2_1 <= AEbuf_2_1_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1446) begin
            mx2_2_2 <= BFbuf_e;
          end else begin
            mx2_2_2 <= AEbuf_2_2_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1559) begin
            mx2_2_3 <= BFbuf_e;
          end else begin
            mx2_2_3 <= AEbuf_2_3_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1672) begin
            mx2_2_4 <= BFbuf_e;
          end else begin
            mx2_2_4 <= AEbuf_2_4_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1785) begin
            mx2_2_5 <= BFbuf_e;
          end else begin
            mx2_2_5 <= AEbuf_2_5_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1898) begin
            mx2_2_6 <= BFbuf_e;
          end else begin
            mx2_2_6 <= AEbuf_2_6_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_2011) begin
            mx2_2_7 <= BFbuf_e;
          end else begin
            mx2_2_7 <= AEbuf_2_7_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1232) begin
            mx2_3_0 <= BFbuf_e;
          end else begin
            mx2_3_0 <= AEbuf_3_0_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1345) begin
            mx2_3_1 <= BFbuf_e;
          end else begin
            mx2_3_1 <= AEbuf_3_1_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1458) begin
            mx2_3_2 <= BFbuf_e;
          end else begin
            mx2_3_2 <= AEbuf_3_2_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1571) begin
            mx2_3_3 <= BFbuf_e;
          end else begin
            mx2_3_3 <= AEbuf_3_3_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1684) begin
            mx2_3_4 <= BFbuf_e;
          end else begin
            mx2_3_4 <= AEbuf_3_4_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1797) begin
            mx2_3_5 <= BFbuf_e;
          end else begin
            mx2_3_5 <= AEbuf_3_5_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1910) begin
            mx2_3_6 <= BFbuf_e;
          end else begin
            mx2_3_6 <= AEbuf_3_6_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_2023) begin
            mx2_3_7 <= BFbuf_e;
          end else begin
            mx2_3_7 <= AEbuf_3_7_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1244) begin
            mx2_4_0 <= BFbuf_e;
          end else begin
            mx2_4_0 <= AEbuf_4_0_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1357) begin
            mx2_4_1 <= BFbuf_e;
          end else begin
            mx2_4_1 <= AEbuf_4_1_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1470) begin
            mx2_4_2 <= BFbuf_e;
          end else begin
            mx2_4_2 <= AEbuf_4_2_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1583) begin
            mx2_4_3 <= BFbuf_e;
          end else begin
            mx2_4_3 <= AEbuf_4_3_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1696) begin
            mx2_4_4 <= BFbuf_e;
          end else begin
            mx2_4_4 <= AEbuf_4_4_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1809) begin
            mx2_4_5 <= BFbuf_e;
          end else begin
            mx2_4_5 <= AEbuf_4_5_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1922) begin
            mx2_4_6 <= BFbuf_e;
          end else begin
            mx2_4_6 <= AEbuf_4_6_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_2035) begin
            mx2_4_7 <= BFbuf_e;
          end else begin
            mx2_4_7 <= AEbuf_4_7_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1256) begin
            mx2_5_0 <= BFbuf_e;
          end else begin
            mx2_5_0 <= AEbuf_5_0_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1369) begin
            mx2_5_1 <= BFbuf_e;
          end else begin
            mx2_5_1 <= AEbuf_5_1_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1482) begin
            mx2_5_2 <= BFbuf_e;
          end else begin
            mx2_5_2 <= AEbuf_5_2_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1595) begin
            mx2_5_3 <= BFbuf_e;
          end else begin
            mx2_5_3 <= AEbuf_5_3_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1708) begin
            mx2_5_4 <= BFbuf_e;
          end else begin
            mx2_5_4 <= AEbuf_5_4_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1821) begin
            mx2_5_5 <= BFbuf_e;
          end else begin
            mx2_5_5 <= AEbuf_5_5_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1934) begin
            mx2_5_6 <= BFbuf_e;
          end else begin
            mx2_5_6 <= AEbuf_5_6_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_2047) begin
            mx2_5_7 <= BFbuf_e;
          end else begin
            mx2_5_7 <= AEbuf_5_7_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1268) begin
            mx2_6_0 <= BFbuf_e;
          end else begin
            mx2_6_0 <= AEbuf_6_0_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1381) begin
            mx2_6_1 <= BFbuf_e;
          end else begin
            mx2_6_1 <= AEbuf_6_1_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1494) begin
            mx2_6_2 <= BFbuf_e;
          end else begin
            mx2_6_2 <= AEbuf_6_2_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1607) begin
            mx2_6_3 <= BFbuf_e;
          end else begin
            mx2_6_3 <= AEbuf_6_3_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1720) begin
            mx2_6_4 <= BFbuf_e;
          end else begin
            mx2_6_4 <= AEbuf_6_4_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1833) begin
            mx2_6_5 <= BFbuf_e;
          end else begin
            mx2_6_5 <= AEbuf_6_5_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1946) begin
            mx2_6_6 <= BFbuf_e;
          end else begin
            mx2_6_6 <= AEbuf_6_6_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_2059) begin
            mx2_6_7 <= BFbuf_e;
          end else begin
            mx2_6_7 <= AEbuf_6_7_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1280) begin
            mx2_7_0 <= BFbuf_e;
          end else begin
            mx2_7_0 <= AEbuf_7_0_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1393) begin
            mx2_7_1 <= BFbuf_e;
          end else begin
            mx2_7_1 <= AEbuf_7_1_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1506) begin
            mx2_7_2 <= BFbuf_e;
          end else begin
            mx2_7_2 <= AEbuf_7_2_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1619) begin
            mx2_7_3 <= BFbuf_e;
          end else begin
            mx2_7_3 <= AEbuf_7_3_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1732) begin
            mx2_7_4 <= BFbuf_e;
          end else begin
            mx2_7_4 <= AEbuf_7_4_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1845) begin
            mx2_7_5 <= BFbuf_e;
          end else begin
            mx2_7_5 <= AEbuf_7_5_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1958) begin
            mx2_7_6 <= BFbuf_e;
          end else begin
            mx2_7_6 <= AEbuf_7_6_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_2071) begin
            mx2_7_7 <= BFbuf_e;
          end else begin
            mx2_7_7 <= AEbuf_7_7_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1200) begin
            ab2_0_0 <= _T_1202;
          end else begin
            ab2_0_0 <= _T_1198;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1313) begin
            ab2_0_1 <= _T_1315;
          end else begin
            ab2_0_1 <= _T_1311;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1426) begin
            ab2_0_2 <= _T_1428;
          end else begin
            ab2_0_2 <= _T_1424;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1539) begin
            ab2_0_3 <= _T_1541;
          end else begin
            ab2_0_3 <= _T_1537;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1652) begin
            ab2_0_4 <= _T_1654;
          end else begin
            ab2_0_4 <= _T_1650;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1765) begin
            ab2_0_5 <= _T_1767;
          end else begin
            ab2_0_5 <= _T_1763;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1878) begin
            ab2_0_6 <= _T_1880;
          end else begin
            ab2_0_6 <= _T_1876;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1991) begin
            ab2_0_7 <= _T_1993;
          end else begin
            ab2_0_7 <= _T_1989;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1212) begin
            ab2_1_0 <= _T_1214;
          end else begin
            ab2_1_0 <= _T_1210;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1325) begin
            ab2_1_1 <= _T_1327;
          end else begin
            ab2_1_1 <= _T_1323;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1438) begin
            ab2_1_2 <= _T_1440;
          end else begin
            ab2_1_2 <= _T_1436;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1551) begin
            ab2_1_3 <= _T_1553;
          end else begin
            ab2_1_3 <= _T_1549;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1664) begin
            ab2_1_4 <= _T_1666;
          end else begin
            ab2_1_4 <= _T_1662;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1777) begin
            ab2_1_5 <= _T_1779;
          end else begin
            ab2_1_5 <= _T_1775;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1890) begin
            ab2_1_6 <= _T_1892;
          end else begin
            ab2_1_6 <= _T_1888;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_2003) begin
            ab2_1_7 <= _T_2005;
          end else begin
            ab2_1_7 <= _T_2001;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1224) begin
            ab2_2_0 <= _T_1226;
          end else begin
            ab2_2_0 <= _T_1222;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1337) begin
            ab2_2_1 <= _T_1339;
          end else begin
            ab2_2_1 <= _T_1335;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1450) begin
            ab2_2_2 <= _T_1452;
          end else begin
            ab2_2_2 <= _T_1448;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1563) begin
            ab2_2_3 <= _T_1565;
          end else begin
            ab2_2_3 <= _T_1561;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1676) begin
            ab2_2_4 <= _T_1678;
          end else begin
            ab2_2_4 <= _T_1674;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1789) begin
            ab2_2_5 <= _T_1791;
          end else begin
            ab2_2_5 <= _T_1787;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1902) begin
            ab2_2_6 <= _T_1904;
          end else begin
            ab2_2_6 <= _T_1900;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_2015) begin
            ab2_2_7 <= _T_2017;
          end else begin
            ab2_2_7 <= _T_2013;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1236) begin
            ab2_3_0 <= _T_1238;
          end else begin
            ab2_3_0 <= _T_1234;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1349) begin
            ab2_3_1 <= _T_1351;
          end else begin
            ab2_3_1 <= _T_1347;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1462) begin
            ab2_3_2 <= _T_1464;
          end else begin
            ab2_3_2 <= _T_1460;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1575) begin
            ab2_3_3 <= _T_1577;
          end else begin
            ab2_3_3 <= _T_1573;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1688) begin
            ab2_3_4 <= _T_1690;
          end else begin
            ab2_3_4 <= _T_1686;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1801) begin
            ab2_3_5 <= _T_1803;
          end else begin
            ab2_3_5 <= _T_1799;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1914) begin
            ab2_3_6 <= _T_1916;
          end else begin
            ab2_3_6 <= _T_1912;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_2027) begin
            ab2_3_7 <= _T_2029;
          end else begin
            ab2_3_7 <= _T_2025;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1248) begin
            ab2_4_0 <= _T_1250;
          end else begin
            ab2_4_0 <= _T_1246;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1361) begin
            ab2_4_1 <= _T_1363;
          end else begin
            ab2_4_1 <= _T_1359;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1474) begin
            ab2_4_2 <= _T_1476;
          end else begin
            ab2_4_2 <= _T_1472;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1587) begin
            ab2_4_3 <= _T_1589;
          end else begin
            ab2_4_3 <= _T_1585;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1700) begin
            ab2_4_4 <= _T_1702;
          end else begin
            ab2_4_4 <= _T_1698;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1813) begin
            ab2_4_5 <= _T_1815;
          end else begin
            ab2_4_5 <= _T_1811;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1926) begin
            ab2_4_6 <= _T_1928;
          end else begin
            ab2_4_6 <= _T_1924;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_2039) begin
            ab2_4_7 <= _T_2041;
          end else begin
            ab2_4_7 <= _T_2037;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1260) begin
            ab2_5_0 <= _T_1262;
          end else begin
            ab2_5_0 <= _T_1258;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1373) begin
            ab2_5_1 <= _T_1375;
          end else begin
            ab2_5_1 <= _T_1371;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1486) begin
            ab2_5_2 <= _T_1488;
          end else begin
            ab2_5_2 <= _T_1484;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1599) begin
            ab2_5_3 <= _T_1601;
          end else begin
            ab2_5_3 <= _T_1597;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1712) begin
            ab2_5_4 <= _T_1714;
          end else begin
            ab2_5_4 <= _T_1710;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1825) begin
            ab2_5_5 <= _T_1827;
          end else begin
            ab2_5_5 <= _T_1823;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1938) begin
            ab2_5_6 <= _T_1940;
          end else begin
            ab2_5_6 <= _T_1936;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_2051) begin
            ab2_5_7 <= _T_2053;
          end else begin
            ab2_5_7 <= _T_2049;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1272) begin
            ab2_6_0 <= _T_1274;
          end else begin
            ab2_6_0 <= _T_1270;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1385) begin
            ab2_6_1 <= _T_1387;
          end else begin
            ab2_6_1 <= _T_1383;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1498) begin
            ab2_6_2 <= _T_1500;
          end else begin
            ab2_6_2 <= _T_1496;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1611) begin
            ab2_6_3 <= _T_1613;
          end else begin
            ab2_6_3 <= _T_1609;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1724) begin
            ab2_6_4 <= _T_1726;
          end else begin
            ab2_6_4 <= _T_1722;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1837) begin
            ab2_6_5 <= _T_1839;
          end else begin
            ab2_6_5 <= _T_1835;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1950) begin
            ab2_6_6 <= _T_1952;
          end else begin
            ab2_6_6 <= _T_1948;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_2063) begin
            ab2_6_7 <= _T_2065;
          end else begin
            ab2_6_7 <= _T_2061;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1284) begin
            ab2_7_0 <= _T_1286;
          end else begin
            ab2_7_0 <= _T_1282;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1397) begin
            ab2_7_1 <= _T_1399;
          end else begin
            ab2_7_1 <= _T_1395;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1510) begin
            ab2_7_2 <= _T_1512;
          end else begin
            ab2_7_2 <= _T_1508;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1623) begin
            ab2_7_3 <= _T_1625;
          end else begin
            ab2_7_3 <= _T_1621;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1736) begin
            ab2_7_4 <= _T_1738;
          end else begin
            ab2_7_4 <= _T_1734;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1849) begin
            ab2_7_5 <= _T_1851;
          end else begin
            ab2_7_5 <= _T_1847;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1962) begin
            ab2_7_6 <= _T_1964;
          end else begin
            ab2_7_6 <= _T_1960;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_2075) begin
            ab2_7_7 <= _T_2077;
          end else begin
            ab2_7_7 <= _T_2073;
          end
        end
      end
    end
    tm8_0_0 <= $signed(_GEN_4987);
    tm8_0_1 <= $signed(_GEN_4988);
    tm8_0_2 <= $signed(_GEN_4989);
    tm8_0_3 <= $signed(_GEN_4990);
    tm8_0_4 <= $signed(_GEN_4991);
    tm8_0_5 <= $signed(_GEN_4992);
    tm8_0_6 <= $signed(_GEN_4993);
    tm8_0_7 <= $signed(_GEN_4994);
    tm8_1_0 <= $signed(_GEN_4995);
    tm8_1_1 <= $signed(_GEN_4996);
    tm8_1_2 <= $signed(_GEN_4997);
    tm8_1_3 <= $signed(_GEN_4998);
    tm8_1_4 <= $signed(_GEN_4999);
    tm8_1_5 <= $signed(_GEN_5000);
    tm8_1_6 <= $signed(_GEN_5001);
    tm8_1_7 <= $signed(_GEN_5002);
    tm8_2_0 <= $signed(_GEN_5003);
    tm8_2_1 <= $signed(_GEN_5004);
    tm8_2_2 <= $signed(_GEN_5005);
    tm8_2_3 <= $signed(_GEN_5006);
    tm8_2_4 <= $signed(_GEN_5007);
    tm8_2_5 <= $signed(_GEN_5008);
    tm8_2_6 <= $signed(_GEN_5009);
    tm8_2_7 <= $signed(_GEN_5010);
    tm8_3_0 <= $signed(_GEN_5011);
    tm8_3_1 <= $signed(_GEN_5012);
    tm8_3_2 <= $signed(_GEN_5013);
    tm8_3_3 <= $signed(_GEN_5014);
    tm8_3_4 <= $signed(_GEN_5015);
    tm8_3_5 <= $signed(_GEN_5016);
    tm8_3_6 <= $signed(_GEN_5017);
    tm8_3_7 <= $signed(_GEN_5018);
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1300) begin
            tm9_0_0 <= tm8_0_0;
          end else begin
            tm9_0_0 <= tm8_1_0;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1413) begin
            tm9_0_1 <= tm8_0_1;
          end else begin
            tm9_0_1 <= tm8_1_1;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1526) begin
            tm9_0_2 <= tm8_0_2;
          end else begin
            tm9_0_2 <= tm8_1_2;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1639) begin
            tm9_0_3 <= tm8_0_3;
          end else begin
            tm9_0_3 <= tm8_1_3;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1752) begin
            tm9_0_4 <= tm8_0_4;
          end else begin
            tm9_0_4 <= tm8_1_4;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1865) begin
            tm9_0_5 <= tm8_0_5;
          end else begin
            tm9_0_5 <= tm8_1_5;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1978) begin
            tm9_0_6 <= tm8_0_6;
          end else begin
            tm9_0_6 <= tm8_1_6;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_2091) begin
            tm9_0_7 <= tm8_0_7;
          end else begin
            tm9_0_7 <= tm8_1_7;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1302) begin
            tm9_1_0 <= tm8_2_0;
          end else begin
            tm9_1_0 <= tm8_3_0;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1415) begin
            tm9_1_1 <= tm8_2_1;
          end else begin
            tm9_1_1 <= tm8_3_1;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1528) begin
            tm9_1_2 <= tm8_2_2;
          end else begin
            tm9_1_2 <= tm8_3_2;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1641) begin
            tm9_1_3 <= tm8_2_3;
          end else begin
            tm9_1_3 <= tm8_3_3;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1754) begin
            tm9_1_4 <= tm8_2_4;
          end else begin
            tm9_1_4 <= tm8_3_4;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1867) begin
            tm9_1_5 <= tm8_2_5;
          end else begin
            tm9_1_5 <= tm8_3_5;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1980) begin
            tm9_1_6 <= tm8_2_6;
          end else begin
            tm9_1_6 <= tm8_3_6;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_2093) begin
            tm9_1_7 <= tm8_2_7;
          end else begin
            tm9_1_7 <= tm8_3_7;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1304) begin
            tma_0_0 <= tm9_0_0;
          end else begin
            tma_0_0 <= tm9_1_0;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1417) begin
            tma_0_1 <= tm9_0_1;
          end else begin
            tma_0_1 <= tm9_1_1;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1530) begin
            tma_0_2 <= tm9_0_2;
          end else begin
            tma_0_2 <= tm9_1_2;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1643) begin
            tma_0_3 <= tm9_0_3;
          end else begin
            tma_0_3 <= tm9_1_3;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1756) begin
            tma_0_4 <= tm9_0_4;
          end else begin
            tma_0_4 <= tm9_1_4;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1869) begin
            tma_0_5 <= tm9_0_5;
          end else begin
            tma_0_5 <= tm9_1_5;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1982) begin
            tma_0_6 <= tm9_0_6;
          end else begin
            tma_0_6 <= tm9_1_6;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_2095) begin
            tma_0_7 <= tm9_0_7;
          end else begin
            tma_0_7 <= tm9_1_7;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          tmb_0_0 <= tma_0_0;
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          tmb_0_1 <= tma_0_1;
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          tmb_0_2 <= tma_0_2;
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          tmb_0_3 <= tma_0_3;
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          tmb_0_4 <= tma_0_4;
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          tmb_0_5 <= tma_0_5;
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          tmb_0_6 <= tma_0_6;
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          tmb_0_7 <= tma_0_7;
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          tmc_0_0 <= tmb_0_0;
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          tmc_0_1 <= tmb_0_1;
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          tmc_0_2 <= tmb_0_2;
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          tmc_0_3 <= tmb_0_3;
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          tmc_0_4 <= tmb_0_4;
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          tmc_0_5 <= tmb_0_5;
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          tmc_0_6 <= tmb_0_6;
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          tmc_0_7 <= tmb_0_7;
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1307) begin
            best_0 <= tmc_0_0;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1420) begin
            best_1 <= tmc_0_1;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1533) begin
            best_2 <= tmc_0_2;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1646) begin
            best_3 <= tmc_0_3;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1759) begin
            best_4 <= tmc_0_4;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1872) begin
            best_5 <= tmc_0_5;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_1985) begin
            best_6 <= tmc_0_6;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_2098) begin
            best_7 <= tmc_0_7;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          bestBufe_0 <= best_0;
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          bestBufe_1 <= best_1;
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          bestBufe_2 <= best_2;
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          bestBufe_3 <= best_3;
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          bestBufe_4 <= best_4;
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          bestBufe_5 <= best_5;
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          bestBufe_6 <= best_6;
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          bestBufe_7 <= best_7;
        end
      end
    end
    if (reset) begin
      r <= 2'h0;
    end else begin
      if (_T_451) begin
        if (_T_452) begin
          if (_T_463) begin
            if (_T_466) begin
              if (_T_2102) begin
                r <= _T_2104;
              end else begin
                r <= 2'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      c <= 2'h0;
    end else begin
      if (_T_451) begin
        if (_T_452) begin
          if (_T_463) begin
            if (_T_466) begin
              if (!(_T_2102)) begin
                if (_T_2105) begin
                  c <= _T_2107;
                end else begin
                  c <= 2'h0;
                end
              end
            end
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_487) begin
            BFbuf_e <= io_lof_bits_e;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_487) begin
            BFbuf_a <= io_lof_bits_a;
          end
        end
      end
    end
    if (reset) begin
      load_i <= 5'h0;
    end else begin
      if (_T_2) begin
        if (io_modeLoad) begin
          if (_T_3) begin
            if (!(lastLoad)) begin
              if (!(_T_398)) begin
                if (_T_401) begin
                  load_i <= _T_403;
                end else begin
                  load_i <= 5'h0;
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      load_j <= 5'h0;
    end else begin
      if (_T_2) begin
        if (io_modeLoad) begin
          if (_T_3) begin
            if (!(lastLoad)) begin
              if (_T_398) begin
                load_j <= _T_400;
              end else begin
                load_j <= 5'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      doneLoading <= 1'h0;
    end else begin
      if (_T_2) begin
        if (io_modeLoad) begin
          if (_T_3) begin
            if (lastLoad) begin
              doneLoading <= 1'h1;
            end
          end
        end else begin
          doneLoading <= 1'h1;
        end
      end
    end
    if (reset) begin
      lastLoad <= 1'h0;
    end else begin
      if (_T_2) begin
        if (io_modeLoad) begin
          if (_T_3) begin
            if (!(lastLoad)) begin
              if (!(_T_398)) begin
                if (!(_T_401)) begin
                  lastLoad <= 1'h1;
                end
              end
            end
          end
        end
      end
    end
    if (_T_2) begin
      if (io_modeLoad) begin
        if (_T_3) begin
          if (!(lastLoad)) begin
            prev_lo_i <= _T_388;
          end
        end
      end
    end
    if (_T_2) begin
      if (io_modeLoad) begin
        if (_T_3) begin
          if (!(lastLoad)) begin
            prev_lo_j <= _T_390;
          end
        end
      end
    end
    if (_T_2) begin
      if (io_modeLoad) begin
        if (_T_3) begin
          if (!(lastLoad)) begin
            prev_idx <= _T_397;
          end
        end
      end
    end
    if (_T_2) begin
      if (io_modeLoad) begin
        if (_T_3) begin
          if (!(lastLoad)) begin
            slcBuf_e <= io_slc_bits_e;
          end
        end
      end
    end
    if (_T_2) begin
      if (io_modeLoad) begin
        if (_T_3) begin
          if (!(lastLoad)) begin
            slcBuf_a <= io_slc_bits_a;
          end
        end
      end
    end
    if (reset) begin
      slcValid <= 1'h0;
    end else begin
      if (_T_2) begin
        if (io_modeLoad) begin
          if (_T_3) begin
            if (!(lastLoad)) begin
              slcValid <= 1'h1;
            end
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_0_0_e <= _T_501;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_0_0_a <= _T_500;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_0_1_e <= _T_589;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_0_1_a <= _T_588;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_0_2_e <= _T_677;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_0_2_a <= _T_676;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_0_3_e <= _T_765;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_0_3_a <= _T_764;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_0_4_e <= _T_853;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_0_4_a <= _T_852;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_0_5_e <= _T_941;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_0_5_a <= _T_940;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_0_6_e <= _T_1029;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_0_6_a <= _T_1028;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_0_7_e <= _T_1117;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_0_7_a <= _T_1116;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_1_0_e <= _T_512;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_1_0_a <= _T_511;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_1_1_e <= _T_600;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_1_1_a <= _T_599;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_1_2_e <= _T_688;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_1_2_a <= _T_687;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_1_3_e <= _T_776;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_1_3_a <= _T_775;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_1_4_e <= _T_864;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_1_4_a <= _T_863;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_1_5_e <= _T_952;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_1_5_a <= _T_951;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_1_6_e <= _T_1040;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_1_6_a <= _T_1039;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_1_7_e <= _T_1128;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_1_7_a <= _T_1127;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_2_0_e <= _T_523;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_2_0_a <= _T_522;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_2_1_e <= _T_611;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_2_1_a <= _T_610;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_2_2_e <= _T_699;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_2_2_a <= _T_698;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_2_3_e <= _T_787;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_2_3_a <= _T_786;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_2_4_e <= _T_875;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_2_4_a <= _T_874;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_2_5_e <= _T_963;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_2_5_a <= _T_962;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_2_6_e <= _T_1051;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_2_6_a <= _T_1050;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_2_7_e <= _T_1139;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_2_7_a <= _T_1138;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_3_0_e <= _T_534;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_3_0_a <= _T_533;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_3_1_e <= _T_622;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_3_1_a <= _T_621;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_3_2_e <= _T_710;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_3_2_a <= _T_709;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_3_3_e <= _T_798;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_3_3_a <= _T_797;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_3_4_e <= _T_886;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_3_4_a <= _T_885;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_3_5_e <= _T_974;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_3_5_a <= _T_973;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_3_6_e <= _T_1062;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_3_6_a <= _T_1061;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_3_7_e <= _T_1150;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_3_7_a <= _T_1149;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_4_0_e <= _T_545;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_4_0_a <= _T_544;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_4_1_e <= _T_633;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_4_1_a <= _T_632;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_4_2_e <= _T_721;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_4_2_a <= _T_720;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_4_3_e <= _T_809;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_4_3_a <= _T_808;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_4_4_e <= _T_897;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_4_4_a <= _T_896;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_4_5_e <= _T_985;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_4_5_a <= _T_984;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_4_6_e <= _T_1073;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_4_6_a <= _T_1072;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_4_7_e <= _T_1161;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_4_7_a <= _T_1160;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_5_0_e <= _T_556;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_5_0_a <= _T_555;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_5_1_e <= _T_644;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_5_1_a <= _T_643;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_5_2_e <= _T_732;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_5_2_a <= _T_731;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_5_3_e <= _T_820;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_5_3_a <= _T_819;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_5_4_e <= _T_908;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_5_4_a <= _T_907;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_5_5_e <= _T_996;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_5_5_a <= _T_995;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_5_6_e <= _T_1084;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_5_6_a <= _T_1083;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_5_7_e <= _T_1172;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_5_7_a <= _T_1171;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_6_0_e <= _T_567;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_6_0_a <= _T_566;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_6_1_e <= _T_655;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_6_1_a <= _T_654;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_6_2_e <= _T_743;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_6_2_a <= _T_742;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_6_3_e <= _T_831;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_6_3_a <= _T_830;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_6_4_e <= _T_919;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_6_4_a <= _T_918;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_6_5_e <= _T_1007;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_6_5_a <= _T_1006;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_6_6_e <= _T_1095;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_6_6_a <= _T_1094;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_6_7_e <= _T_1183;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_6_7_a <= _T_1182;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_7_0_e <= _T_578;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_7_0_a <= _T_577;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_7_1_e <= _T_666;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_7_1_a <= _T_665;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_7_2_e <= _T_754;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_7_2_a <= _T_753;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_7_3_e <= _T_842;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_7_3_a <= _T_841;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_7_4_e <= _T_930;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_7_4_a <= _T_929;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_7_5_e <= _T_1018;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_7_5_a <= _T_1017;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_7_6_e <= _T_1106;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_7_6_a <= _T_1105;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_7_7_e <= _T_1194;
          end
        end
      end
    end
    if (_T_451) begin
      if (_T_452) begin
        if (_T_463) begin
          if (_T_466) begin
            AEbuf_7_7_a <= _T_1193;
          end
        end
      end
    end
    if (reset) begin
      _T_405 <= 1'h0;
    end else begin
      if (_T_451) begin
        if (_T_452) begin
          if (_T_463) begin
            _T_405 <= _T_466;
          end
        end
      end
    end
    if (reset) begin
      _T_406 <= 1'h0;
    end else begin
      if (_T_451) begin
        if (_T_452) begin
          if (_T_463) begin
            _T_406 <= _T_405;
          end
        end
      end
    end
    if (reset) begin
      _T_407 <= 1'h0;
    end else begin
      if (_T_451) begin
        if (_T_452) begin
          if (_T_463) begin
            _T_407 <= _T_406;
          end
        end
      end
    end
    if (reset) begin
      _T_408 <= 1'h0;
    end else begin
      if (_T_451) begin
        if (_T_452) begin
          if (_T_463) begin
            _T_408 <= _T_407;
          end
        end
      end
    end
    if (reset) begin
      _T_409 <= 1'h0;
    end else begin
      if (_T_451) begin
        if (_T_452) begin
          if (_T_463) begin
            _T_409 <= _T_408;
          end
        end
      end
    end
    if (reset) begin
      _T_410 <= 1'h0;
    end else begin
      if (_T_451) begin
        if (_T_452) begin
          if (_T_463) begin
            _T_410 <= _T_409;
          end
        end
      end
    end
    if (reset) begin
      _T_411 <= 1'h0;
    end else begin
      if (_T_451) begin
        if (_T_452) begin
          if (_T_463) begin
            _T_411 <= _T_410;
          end
        end
      end
    end
    if (reset) begin
      _T_412 <= 1'h0;
    end else begin
      if (_T_451) begin
        if (_T_452) begin
          if (_T_463) begin
            _T_412 <= _T_411;
          end
        end
      end
    end
    if (reset) begin
      _T_413 <= 1'h0;
    end else begin
      if (_T_451) begin
        if (_T_452) begin
          if (_T_463) begin
            _T_413 <= _T_412;
          end
        end
      end
    end
    if (reset) begin
      _T_414 <= 1'h0;
    end else begin
      if (_T_451) begin
        if (_T_452) begin
          if (_T_463) begin
            _T_414 <= _T_413;
          end
        end
      end
    end
    if (reset) begin
      _T_415 <= 1'h0;
    end else begin
      if (_T_451) begin
        if (_T_452) begin
          if (_T_463) begin
            _T_415 <= _T_414;
          end
        end
      end
    end
    if (reset) begin
      _T_416 <= 1'h0;
    end else begin
      if (_T_451) begin
        if (_T_452) begin
          if (_T_463) begin
            _T_416 <= _T_415;
          end
        end
      end
    end
    if (reset) begin
      _T_417 <= 1'h0;
    end else begin
      if (_T_451) begin
        if (_T_452) begin
          if (_T_463) begin
            _T_417 <= _T_416;
          end
        end
      end
    end
    if (reset) begin
      _T_418 <= 1'h0;
    end else begin
      if (_T_451) begin
        if (_T_452) begin
          if (_T_463) begin
            _T_418 <= _T_417;
          end
        end
      end
    end
    if (reset) begin
      _T_421 <= 1'h0;
    end else begin
      if (_T_451) begin
        if (_T_452) begin
          if (_T_463) begin
            _T_421 <= _T_471;
          end
        end
      end
    end
    if (reset) begin
      _T_422 <= 1'h0;
    end else begin
      if (_T_451) begin
        if (_T_452) begin
          if (_T_463) begin
            _T_422 <= _T_421;
          end
        end
      end
    end
    if (reset) begin
      _T_423 <= 1'h0;
    end else begin
      if (_T_451) begin
        if (_T_452) begin
          if (_T_463) begin
            _T_423 <= _T_422;
          end
        end
      end
    end
    if (reset) begin
      _T_424 <= 1'h0;
    end else begin
      if (_T_451) begin
        if (_T_452) begin
          if (_T_463) begin
            _T_424 <= _T_423;
          end
        end
      end
    end
    if (reset) begin
      _T_425 <= 1'h0;
    end else begin
      if (_T_451) begin
        if (_T_452) begin
          if (_T_463) begin
            _T_425 <= _T_424;
          end
        end
      end
    end
    if (reset) begin
      _T_426 <= 1'h0;
    end else begin
      if (_T_451) begin
        if (_T_452) begin
          if (_T_463) begin
            _T_426 <= _T_425;
          end
        end
      end
    end
    if (reset) begin
      _T_427 <= 1'h0;
    end else begin
      if (_T_451) begin
        if (_T_452) begin
          if (_T_463) begin
            _T_427 <= _T_426;
          end
        end
      end
    end
    if (reset) begin
      _T_428 <= 1'h0;
    end else begin
      if (_T_451) begin
        if (_T_452) begin
          if (_T_463) begin
            _T_428 <= _T_427;
          end
        end
      end
    end
    if (reset) begin
      _T_429 <= 1'h0;
    end else begin
      if (_T_451) begin
        if (_T_452) begin
          if (_T_463) begin
            _T_429 <= _T_428;
          end
        end
      end
    end
    if (reset) begin
      _T_430 <= 1'h0;
    end else begin
      if (_T_451) begin
        if (_T_452) begin
          if (_T_463) begin
            _T_430 <= _T_429;
          end
        end
      end
    end
    if (reset) begin
      _T_431 <= 1'h0;
    end else begin
      if (_T_451) begin
        if (_T_452) begin
          if (_T_463) begin
            _T_431 <= _T_430;
          end
        end
      end
    end
    if (reset) begin
      _T_432 <= 1'h0;
    end else begin
      if (_T_451) begin
        if (_T_452) begin
          if (_T_463) begin
            _T_432 <= _T_431;
          end
        end
      end
    end
    if (reset) begin
      _T_433 <= 1'h0;
    end else begin
      if (_T_451) begin
        if (_T_452) begin
          if (_T_463) begin
            _T_433 <= _T_432;
          end
        end
      end
    end
    if (reset) begin
      _T_434 <= 1'h0;
    end else begin
      if (_T_451) begin
        if (_T_452) begin
          if (_T_463) begin
            _T_434 <= _T_433;
          end
        end
      end
    end
    if (reset) begin
      _T_437 <= 1'h0;
    end else begin
      if (_T_451) begin
        if (_T_452) begin
          if (_T_463) begin
            _T_437 <= _T_476;
          end
        end
      end
    end
    if (reset) begin
      _T_438 <= 1'h0;
    end else begin
      if (_T_451) begin
        if (_T_452) begin
          if (_T_463) begin
            _T_438 <= _T_437;
          end
        end
      end
    end
    if (reset) begin
      _T_439 <= 1'h0;
    end else begin
      if (_T_451) begin
        if (_T_452) begin
          if (_T_463) begin
            _T_439 <= _T_438;
          end
        end
      end
    end
    if (reset) begin
      _T_440 <= 1'h0;
    end else begin
      if (_T_451) begin
        if (_T_452) begin
          if (_T_463) begin
            _T_440 <= _T_439;
          end
        end
      end
    end
    if (reset) begin
      _T_441 <= 1'h0;
    end else begin
      if (_T_451) begin
        if (_T_452) begin
          if (_T_463) begin
            _T_441 <= _T_440;
          end
        end
      end
    end
    if (reset) begin
      _T_442 <= 1'h0;
    end else begin
      if (_T_451) begin
        if (_T_452) begin
          if (_T_463) begin
            _T_442 <= _T_441;
          end
        end
      end
    end
    if (reset) begin
      _T_443 <= 1'h0;
    end else begin
      if (_T_451) begin
        if (_T_452) begin
          if (_T_463) begin
            _T_443 <= _T_442;
          end
        end
      end
    end
    if (reset) begin
      _T_444 <= 1'h0;
    end else begin
      if (_T_451) begin
        if (_T_452) begin
          if (_T_463) begin
            _T_444 <= _T_443;
          end
        end
      end
    end
    if (reset) begin
      _T_445 <= 1'h0;
    end else begin
      if (_T_451) begin
        if (_T_452) begin
          if (_T_463) begin
            _T_445 <= _T_444;
          end
        end
      end
    end
    if (reset) begin
      _T_446 <= 1'h0;
    end else begin
      if (_T_451) begin
        if (_T_452) begin
          if (_T_463) begin
            _T_446 <= _T_445;
          end
        end
      end
    end
    if (reset) begin
      _T_447 <= 1'h0;
    end else begin
      if (_T_451) begin
        if (_T_452) begin
          if (_T_463) begin
            _T_447 <= _T_446;
          end
        end
      end
    end
    if (reset) begin
      _T_448 <= 1'h0;
    end else begin
      if (_T_451) begin
        if (_T_452) begin
          if (_T_463) begin
            _T_448 <= _T_447;
          end
        end
      end
    end
  end
endmodule
module SplitOut(
  input         io_start,
  output        io_out_ready,
  input         io_out_valid,
  input  [15:0] io_out_bits_0,
  input  [15:0] io_out_bits_1,
  input  [15:0] io_out_bits_2,
  input  [15:0] io_out_bits_3,
  input  [15:0] io_out_bits_4,
  input  [15:0] io_out_bits_5,
  input  [15:0] io_out_bits_6,
  input  [15:0] io_out_bits_7,
  input         io_out0_ready,
  output        io_out0_valid,
  output [15:0] io_out0_bits_0,
  output [15:0] io_out0_bits_1,
  output [15:0] io_out0_bits_2,
  output [15:0] io_out0_bits_3,
  output [15:0] io_out0_bits_4,
  output [15:0] io_out0_bits_5,
  output [15:0] io_out0_bits_6,
  output [15:0] io_out0_bits_7,
  input         io_out1_ready,
  output        io_out1_valid,
  output [15:0] io_out1_bits_0,
  output [15:0] io_out1_bits_1,
  output [15:0] io_out1_bits_2,
  output [15:0] io_out1_bits_3,
  output [15:0] io_out1_bits_4,
  output [15:0] io_out1_bits_5,
  output [15:0] io_out1_bits_6,
  output [15:0] io_out1_bits_7
);
  wire  _T; // @[Clamper.scala 23:25]
  wire  _T_1; // @[Clamper.scala 23:42]
  assign _T = io_out_valid & io_out0_ready; // @[Clamper.scala 23:25]
  assign _T_1 = _T & io_out1_ready; // @[Clamper.scala 23:42]
  assign io_out_ready = io_start ? _T_1 : 1'h0; // @[Decoupled.scala 69:20 Clamper.scala 24:20]
  assign io_out0_valid = io_start ? _T_1 : 1'h0; // @[Decoupled.scala 53:20 Clamper.scala 25:21]
  assign io_out0_bits_0 = io_out_bits_0; // @[Clamper.scala 27:20]
  assign io_out0_bits_1 = io_out_bits_1; // @[Clamper.scala 27:20]
  assign io_out0_bits_2 = io_out_bits_2; // @[Clamper.scala 27:20]
  assign io_out0_bits_3 = io_out_bits_3; // @[Clamper.scala 27:20]
  assign io_out0_bits_4 = io_out_bits_4; // @[Clamper.scala 27:20]
  assign io_out0_bits_5 = io_out_bits_5; // @[Clamper.scala 27:20]
  assign io_out0_bits_6 = io_out_bits_6; // @[Clamper.scala 27:20]
  assign io_out0_bits_7 = io_out_bits_7; // @[Clamper.scala 27:20]
  assign io_out1_valid = io_start ? _T_1 : 1'h0; // @[Decoupled.scala 53:20 Clamper.scala 26:21]
  assign io_out1_bits_0 = io_out_bits_0; // @[Clamper.scala 28:20]
  assign io_out1_bits_1 = io_out_bits_1; // @[Clamper.scala 28:20]
  assign io_out1_bits_2 = io_out_bits_2; // @[Clamper.scala 28:20]
  assign io_out1_bits_3 = io_out_bits_3; // @[Clamper.scala 28:20]
  assign io_out1_bits_4 = io_out_bits_4; // @[Clamper.scala 28:20]
  assign io_out1_bits_5 = io_out_bits_5; // @[Clamper.scala 28:20]
  assign io_out1_bits_6 = io_out_bits_6; // @[Clamper.scala 28:20]
  assign io_out1_bits_7 = io_out_bits_7; // @[Clamper.scala 28:20]
endmodule
module ComputeBest(
  input         clock,
  input         reset,
  input         io_start,
  output        io_out0_ready,
  input         io_out0_valid,
  input  [15:0] io_out0_bits_0,
  input  [15:0] io_out0_bits_1,
  input  [15:0] io_out0_bits_2,
  input  [15:0] io_out0_bits_3,
  input  [15:0] io_out0_bits_4,
  input  [15:0] io_out0_bits_5,
  input  [15:0] io_out0_bits_6,
  input  [15:0] io_out0_bits_7,
  input         io_obest_ready,
  output        io_obest_valid,
  output [15:0] io_obest_bits
);
  reg [1:0] jj; // @[Clamper.scala 42:19]
  reg [31:0] _RAND_0;
  reg [15:0] best; // @[Clamper.scala 43:17]
  reg [31:0] _RAND_1;
  reg  validPipe0; // @[Clamper.scala 63:27]
  reg [31:0] _RAND_2;
  reg [1:0] prev_jj0; // @[Clamper.scala 64:25]
  reg [31:0] _RAND_3;
  reg [15:0] m0_0; // @[Clamper.scala 65:15]
  reg [31:0] _RAND_4;
  reg [15:0] m0_1; // @[Clamper.scala 65:15]
  reg [31:0] _RAND_5;
  reg [15:0] m0_2; // @[Clamper.scala 65:15]
  reg [31:0] _RAND_6;
  reg [15:0] m0_3; // @[Clamper.scala 65:15]
  reg [31:0] _RAND_7;
  reg  validPipe1; // @[Clamper.scala 67:27]
  reg [31:0] _RAND_8;
  reg [1:0] prev_jj1; // @[Clamper.scala 68:25]
  reg [31:0] _RAND_9;
  reg [15:0] m1_0; // @[Clamper.scala 69:15]
  reg [31:0] _RAND_10;
  reg [15:0] m1_1; // @[Clamper.scala 69:15]
  reg [31:0] _RAND_11;
  wire  _T_1; // @[Clamper.scala 90:37]
  wire  _T_2; // @[Clamper.scala 90:58]
  wire  _T_3; // @[Clamper.scala 90:23]
  wire  _T_5; // @[Clamper.scala 73:22]
  wire [15:0] _GEN_0; // @[Clamper.scala 73:27]
  wire  _T_7; // @[Clamper.scala 95:53]
  wire  _T_9; // @[Clamper.scala 73:22]
  wire  _T_10; // @[Clamper.scala 73:17]
  wire  _T_11; // @[Clamper.scala 100:23]
  wire  _GEN_5; // @[Clamper.scala 90:78]
  wire  _GEN_7; // @[Clamper.scala 90:78]
  wire  _T_13; // @[Clamper.scala 110:26]
  wire  _T_14; // @[Clamper.scala 110:23]
  wire  _T_16; // @[Clamper.scala 73:22]
  wire  _T_19; // @[Clamper.scala 73:22]
  wire  _GEN_14; // @[Clamper.scala 110:43]
  wire  _T_21; // @[Clamper.scala 129:29]
  wire  _T_22; // @[Clamper.scala 129:26]
  wire  _T_24; // @[Clamper.scala 73:22]
  wire  _T_27; // @[Clamper.scala 73:22]
  wire  _T_30; // @[Clamper.scala 73:22]
  wire  _T_33; // @[Clamper.scala 73:22]
  wire  _T_35; // @[Clamper.scala 145:17]
  wire [1:0] _T_37; // @[Clamper.scala 146:18]
  assign _T_1 = prev_jj1 != 2'h2; // @[Clamper.scala 90:37]
  assign _T_2 = _T_1 | io_obest_ready; // @[Clamper.scala 90:58]
  assign _T_3 = validPipe1 & _T_2; // @[Clamper.scala 90:23]
  assign _T_5 = $signed(m1_0) < $signed(m1_1); // @[Clamper.scala 73:22]
  assign _GEN_0 = _T_5 ? $signed(m1_0) : $signed(m1_1); // @[Clamper.scala 73:27]
  assign _T_7 = prev_jj1 == 2'h0; // @[Clamper.scala 95:53]
  assign _T_9 = $signed(_GEN_0) < $signed(best); // @[Clamper.scala 73:22]
  assign _T_10 = _T_7 | _T_9; // @[Clamper.scala 73:17]
  assign _T_11 = prev_jj1 == 2'h2; // @[Clamper.scala 100:23]
  assign _GEN_5 = _T_3 ? _T_11 : 1'h0; // @[Clamper.scala 90:78]
  assign _GEN_7 = _T_3 ? 1'h0 : validPipe1; // @[Clamper.scala 90:78]
  assign _T_13 = _GEN_7 == 1'h0; // @[Clamper.scala 110:26]
  assign _T_14 = validPipe0 & _T_13; // @[Clamper.scala 110:23]
  assign _T_16 = $signed(m0_0) < $signed(m0_1); // @[Clamper.scala 73:22]
  assign _T_19 = $signed(m0_2) < $signed(m0_3); // @[Clamper.scala 73:22]
  assign _GEN_14 = _T_14 ? 1'h0 : validPipe0; // @[Clamper.scala 110:43]
  assign _T_21 = _GEN_14 == 1'h0; // @[Clamper.scala 129:29]
  assign _T_22 = io_out0_valid & _T_21; // @[Clamper.scala 129:26]
  assign _T_24 = $signed(io_out0_bits_0) < $signed(io_out0_bits_1); // @[Clamper.scala 73:22]
  assign _T_27 = $signed(io_out0_bits_2) < $signed(io_out0_bits_3); // @[Clamper.scala 73:22]
  assign _T_30 = $signed(io_out0_bits_4) < $signed(io_out0_bits_5); // @[Clamper.scala 73:22]
  assign _T_33 = $signed(io_out0_bits_6) < $signed(io_out0_bits_7); // @[Clamper.scala 73:22]
  assign _T_35 = jj != 2'h2; // @[Clamper.scala 145:17]
  assign _T_37 = jj + 2'h1; // @[Clamper.scala 146:18]
  assign io_out0_ready = io_start ? _T_22 : 1'h0; // @[Decoupled.scala 69:20 Clamper.scala 130:21]
  assign io_obest_valid = io_start ? _GEN_5 : 1'h0; // @[Decoupled.scala 53:20 Clamper.scala 101:24]
  assign io_obest_bits = _T_10 ? $signed(_GEN_0) : $signed(best); // @[Clamper.scala 102:23]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  jj = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  best = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  validPipe0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  prev_jj0 = _RAND_3[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  m0_0 = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  m0_1 = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  m0_2 = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  m0_3 = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  validPipe1 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  prev_jj1 = _RAND_9[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  m1_0 = _RAND_10[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  m1_1 = _RAND_11[15:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      jj <= 2'h0;
    end else begin
      if (io_start) begin
        if (_T_22) begin
          if (_T_35) begin
            jj <= _T_37;
          end else begin
            jj <= 2'h0;
          end
        end
      end
    end
    if (io_start) begin
      if (_T_3) begin
        if (_T_10) begin
          if (_T_5) begin
            best <= m1_0;
          end else begin
            best <= m1_1;
          end
        end
      end
    end
    if (reset) begin
      validPipe0 <= 1'h0;
    end else begin
      if (io_start) begin
        if (_T_22) begin
          validPipe0 <= 1'h1;
        end else begin
          if (_T_14) begin
            validPipe0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      prev_jj0 <= 2'h0;
    end else begin
      if (io_start) begin
        if (_T_22) begin
          prev_jj0 <= jj;
        end
      end
    end
    if (io_start) begin
      if (_T_22) begin
        if (_T_24) begin
          m0_0 <= io_out0_bits_0;
        end else begin
          m0_0 <= io_out0_bits_1;
        end
      end
    end
    if (io_start) begin
      if (_T_22) begin
        if (_T_27) begin
          m0_1 <= io_out0_bits_2;
        end else begin
          m0_1 <= io_out0_bits_3;
        end
      end
    end
    if (io_start) begin
      if (_T_22) begin
        if (_T_30) begin
          m0_2 <= io_out0_bits_4;
        end else begin
          m0_2 <= io_out0_bits_5;
        end
      end
    end
    if (io_start) begin
      if (_T_22) begin
        if (_T_33) begin
          m0_3 <= io_out0_bits_6;
        end else begin
          m0_3 <= io_out0_bits_7;
        end
      end
    end
    if (reset) begin
      validPipe1 <= 1'h0;
    end else begin
      if (io_start) begin
        if (_T_14) begin
          validPipe1 <= 1'h1;
        end else begin
          if (_T_3) begin
            validPipe1 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      prev_jj1 <= 2'h0;
    end else begin
      if (io_start) begin
        if (_T_14) begin
          prev_jj1 <= prev_jj0;
        end
      end
    end
    if (io_start) begin
      if (_T_14) begin
        if (_T_16) begin
          m1_0 <= m0_0;
        end else begin
          m1_0 <= m0_1;
        end
      end
    end
    if (io_start) begin
      if (_T_14) begin
        if (_T_19) begin
          m1_1 <= m0_2;
        end else begin
          m1_1 <= m0_3;
        end
      end
    end
  end
endmodule
module SubtractOut(
  input         clock,
  input         reset,
  input         io_start,
  output        io_out1_ready,
  input         io_out1_valid,
  input  [15:0] io_out1_bits_0,
  input  [15:0] io_out1_bits_1,
  input  [15:0] io_out1_bits_2,
  input  [15:0] io_out1_bits_3,
  input  [15:0] io_out1_bits_4,
  input  [15:0] io_out1_bits_5,
  input  [15:0] io_out1_bits_6,
  input  [15:0] io_out1_bits_7,
  output        io_obest_ready,
  input         io_obest_valid,
  input  [15:0] io_obest_bits,
  input         io_res_ready,
  output        io_res_valid,
  output [15:0] io_res_bits_0,
  output [15:0] io_res_bits_1,
  output [15:0] io_res_bits_2,
  output [15:0] io_res_bits_3,
  output [15:0] io_res_bits_4,
  output [15:0] io_res_bits_5,
  output [15:0] io_res_bits_6,
  output [15:0] io_res_bits_7
);
  reg [1:0] jj; // @[Clamper.scala 166:19]
  reg [31:0] _RAND_0;
  reg [15:0] best; // @[Clamper.scala 168:17]
  reg [31:0] _RAND_1;
  wire  _T; // @[Clamper.scala 178:17]
  wire  _T_1; // @[Clamper.scala 178:25]
  wire  _T_2; // @[Clamper.scala 178:44]
  wire  _T_3; // @[Clamper.scala 178:61]
  wire  _T_5; // @[Clamper.scala 180:16]
  wire [15:0] _GEN_1; // @[Clamper.scala 180:25]
  wire [15:0] _T_7; // @[Clamper.scala 188:44]
  wire [15:0] _T_8; // @[Clamper.scala 188:44]
  wire [15:0] _T_11; // @[Clamper.scala 188:44]
  wire [15:0] _T_12; // @[Clamper.scala 188:44]
  wire [15:0] _T_15; // @[Clamper.scala 188:44]
  wire [15:0] _T_16; // @[Clamper.scala 188:44]
  wire [15:0] _T_19; // @[Clamper.scala 188:44]
  wire [15:0] _T_20; // @[Clamper.scala 188:44]
  wire [15:0] _T_23; // @[Clamper.scala 188:44]
  wire [15:0] _T_24; // @[Clamper.scala 188:44]
  wire [15:0] _T_27; // @[Clamper.scala 188:44]
  wire [15:0] _T_28; // @[Clamper.scala 188:44]
  wire [15:0] _T_31; // @[Clamper.scala 188:44]
  wire [15:0] _T_32; // @[Clamper.scala 188:44]
  wire [15:0] _T_35; // @[Clamper.scala 188:44]
  wire [15:0] _T_36; // @[Clamper.scala 188:44]
  wire  _T_38; // @[Clamper.scala 190:17]
  wire [1:0] _T_40; // @[Clamper.scala 191:18]
  wire  _GEN_3; // @[Clamper.scala 178:78]
  assign _T = jj != 2'h0; // @[Clamper.scala 178:17]
  assign _T_1 = _T | io_obest_valid; // @[Clamper.scala 178:25]
  assign _T_2 = _T_1 & io_out1_valid; // @[Clamper.scala 178:44]
  assign _T_3 = _T_2 & io_res_ready; // @[Clamper.scala 178:61]
  assign _T_5 = jj == 2'h0; // @[Clamper.scala 180:16]
  assign _GEN_1 = _T_5 ? $signed(io_obest_bits) : $signed(best); // @[Clamper.scala 180:25]
  assign _T_7 = $signed(io_out1_bits_0) - $signed(_GEN_1); // @[Clamper.scala 188:44]
  assign _T_8 = $signed(_T_7); // @[Clamper.scala 188:44]
  assign _T_11 = $signed(io_out1_bits_1) - $signed(_GEN_1); // @[Clamper.scala 188:44]
  assign _T_12 = $signed(_T_11); // @[Clamper.scala 188:44]
  assign _T_15 = $signed(io_out1_bits_2) - $signed(_GEN_1); // @[Clamper.scala 188:44]
  assign _T_16 = $signed(_T_15); // @[Clamper.scala 188:44]
  assign _T_19 = $signed(io_out1_bits_3) - $signed(_GEN_1); // @[Clamper.scala 188:44]
  assign _T_20 = $signed(_T_19); // @[Clamper.scala 188:44]
  assign _T_23 = $signed(io_out1_bits_4) - $signed(_GEN_1); // @[Clamper.scala 188:44]
  assign _T_24 = $signed(_T_23); // @[Clamper.scala 188:44]
  assign _T_27 = $signed(io_out1_bits_5) - $signed(_GEN_1); // @[Clamper.scala 188:44]
  assign _T_28 = $signed(_T_27); // @[Clamper.scala 188:44]
  assign _T_31 = $signed(io_out1_bits_6) - $signed(_GEN_1); // @[Clamper.scala 188:44]
  assign _T_32 = $signed(_T_31); // @[Clamper.scala 188:44]
  assign _T_35 = $signed(io_out1_bits_7) - $signed(_GEN_1); // @[Clamper.scala 188:44]
  assign _T_36 = $signed(_T_35); // @[Clamper.scala 188:44]
  assign _T_38 = jj != 2'h2; // @[Clamper.scala 190:17]
  assign _T_40 = jj + 2'h1; // @[Clamper.scala 191:18]
  assign _GEN_3 = _T_3 ? _T_5 : 1'h0; // @[Clamper.scala 178:78]
  assign io_out1_ready = io_start ? _T_3 : 1'h0; // @[Decoupled.scala 69:20 Clamper.scala 185:21]
  assign io_obest_ready = io_start ? _GEN_3 : 1'h0; // @[Decoupled.scala 69:20 Clamper.scala 181:24]
  assign io_res_valid = io_start ? _T_3 : 1'h0; // @[Decoupled.scala 53:20 Clamper.scala 186:20]
  assign io_res_bits_0 = $unsigned(_T_8); // @[Clamper.scala 188:24]
  assign io_res_bits_1 = $unsigned(_T_12); // @[Clamper.scala 188:24]
  assign io_res_bits_2 = $unsigned(_T_16); // @[Clamper.scala 188:24]
  assign io_res_bits_3 = $unsigned(_T_20); // @[Clamper.scala 188:24]
  assign io_res_bits_4 = $unsigned(_T_24); // @[Clamper.scala 188:24]
  assign io_res_bits_5 = $unsigned(_T_28); // @[Clamper.scala 188:24]
  assign io_res_bits_6 = $unsigned(_T_32); // @[Clamper.scala 188:24]
  assign io_res_bits_7 = $unsigned(_T_36); // @[Clamper.scala 188:24]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  jj = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  best = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      jj <= 2'h0;
    end else begin
      if (io_start) begin
        if (_T_3) begin
          if (_T_38) begin
            jj <= _T_40;
          end else begin
            jj <= 2'h0;
          end
        end
      end
    end
    if (io_start) begin
      if (_T_3) begin
        if (_T_5) begin
          best <= io_obest_bits;
        end
      end
    end
  end
endmodule
module DecoupledStage(
  input         clock,
  input         reset,
  output        io_inp_ready,
  input         io_inp_valid,
  input  [15:0] io_inp_bits_0,
  input  [15:0] io_inp_bits_1,
  input  [15:0] io_inp_bits_2,
  input  [15:0] io_inp_bits_3,
  input  [15:0] io_inp_bits_4,
  input  [15:0] io_inp_bits_5,
  input  [15:0] io_inp_bits_6,
  input  [15:0] io_inp_bits_7,
  input         io_out_ready,
  output        io_out_valid,
  output [15:0] io_out_bits_0,
  output [15:0] io_out_bits_1,
  output [15:0] io_out_bits_2,
  output [15:0] io_out_bits_3,
  output [15:0] io_out_bits_4,
  output [15:0] io_out_bits_5,
  output [15:0] io_out_bits_6,
  output [15:0] io_out_bits_7
);
  reg  out_valid; // @[DecoupledStage.scala 14:22]
  reg [31:0] _RAND_0;
  reg [15:0] out_bits_0; // @[DecoupledStage.scala 15:21]
  reg [31:0] _RAND_1;
  reg [15:0] out_bits_1; // @[DecoupledStage.scala 15:21]
  reg [31:0] _RAND_2;
  reg [15:0] out_bits_2; // @[DecoupledStage.scala 15:21]
  reg [31:0] _RAND_3;
  reg [15:0] out_bits_3; // @[DecoupledStage.scala 15:21]
  reg [31:0] _RAND_4;
  reg [15:0] out_bits_4; // @[DecoupledStage.scala 15:21]
  reg [31:0] _RAND_5;
  reg [15:0] out_bits_5; // @[DecoupledStage.scala 15:21]
  reg [31:0] _RAND_6;
  reg [15:0] out_bits_6; // @[DecoupledStage.scala 15:21]
  reg [31:0] _RAND_7;
  reg [15:0] out_bits_7; // @[DecoupledStage.scala 15:21]
  reg [31:0] _RAND_8;
  wire  _T; // @[DecoupledStage.scala 20:34]
  wire  _T_2; // @[DecoupledStage.scala 22:31]
  wire  _T_3; // @[DecoupledStage.scala 22:29]
  assign _T = ~ io_out_valid; // @[DecoupledStage.scala 20:34]
  assign _T_2 = ~ io_inp_ready; // @[DecoupledStage.scala 22:31]
  assign _T_3 = io_inp_valid | _T_2; // @[DecoupledStage.scala 22:29]
  assign io_inp_ready = io_out_ready | _T; // @[DecoupledStage.scala 20:16]
  assign io_out_valid = out_valid; // @[DecoupledStage.scala 17:16]
  assign io_out_bits_0 = out_bits_0; // @[DecoupledStage.scala 18:16]
  assign io_out_bits_1 = out_bits_1; // @[DecoupledStage.scala 18:16]
  assign io_out_bits_2 = out_bits_2; // @[DecoupledStage.scala 18:16]
  assign io_out_bits_3 = out_bits_3; // @[DecoupledStage.scala 18:16]
  assign io_out_bits_4 = out_bits_4; // @[DecoupledStage.scala 18:16]
  assign io_out_bits_5 = out_bits_5; // @[DecoupledStage.scala 18:16]
  assign io_out_bits_6 = out_bits_6; // @[DecoupledStage.scala 18:16]
  assign io_out_bits_7 = out_bits_7; // @[DecoupledStage.scala 18:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  out_valid = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  out_bits_0 = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  out_bits_1 = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_bits_2 = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_bits_3 = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  out_bits_4 = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  out_bits_5 = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  out_bits_6 = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  out_bits_7 = _RAND_8[15:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      out_valid <= 1'h0;
    end else begin
      out_valid <= _T_3;
    end
    if (io_inp_ready) begin
      out_bits_0 <= io_inp_bits_0;
    end
    if (io_inp_ready) begin
      out_bits_1 <= io_inp_bits_1;
    end
    if (io_inp_ready) begin
      out_bits_2 <= io_inp_bits_2;
    end
    if (io_inp_ready) begin
      out_bits_3 <= io_inp_bits_3;
    end
    if (io_inp_ready) begin
      out_bits_4 <= io_inp_bits_4;
    end
    if (io_inp_ready) begin
      out_bits_5 <= io_inp_bits_5;
    end
    if (io_inp_ready) begin
      out_bits_6 <= io_inp_bits_6;
    end
    if (io_inp_ready) begin
      out_bits_7 <= io_inp_bits_7;
    end
  end
endmodule
module DecoupledStage_1(
  input         clock,
  input         reset,
  output        io_inp_ready,
  input         io_inp_valid,
  input  [15:0] io_inp_bits,
  input         io_out_ready,
  output        io_out_valid,
  output [15:0] io_out_bits
);
  reg  out_valid; // @[DecoupledStage.scala 14:22]
  reg [31:0] _RAND_0;
  reg [15:0] out_bits; // @[DecoupledStage.scala 15:21]
  reg [31:0] _RAND_1;
  wire  _T; // @[DecoupledStage.scala 20:34]
  wire  _T_2; // @[DecoupledStage.scala 22:31]
  wire  _T_3; // @[DecoupledStage.scala 22:29]
  assign _T = ~ io_out_valid; // @[DecoupledStage.scala 20:34]
  assign _T_2 = ~ io_inp_ready; // @[DecoupledStage.scala 22:31]
  assign _T_3 = io_inp_valid | _T_2; // @[DecoupledStage.scala 22:29]
  assign io_inp_ready = io_out_ready | _T; // @[DecoupledStage.scala 20:16]
  assign io_out_valid = out_valid; // @[DecoupledStage.scala 17:16]
  assign io_out_bits = out_bits; // @[DecoupledStage.scala 18:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  out_valid = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  out_bits = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      out_valid <= 1'h0;
    end else begin
      out_valid <= _T_3;
    end
    if (io_inp_ready) begin
      out_bits <= io_inp_bits;
    end
  end
endmodule
module Queue(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [15:0] io_enq_bits_0,
  input  [15:0] io_enq_bits_1,
  input  [15:0] io_enq_bits_2,
  input  [15:0] io_enq_bits_3,
  input  [15:0] io_enq_bits_4,
  input  [15:0] io_enq_bits_5,
  input  [15:0] io_enq_bits_6,
  input  [15:0] io_enq_bits_7,
  input         io_deq_ready,
  output        io_deq_valid,
  output [15:0] io_deq_bits_0,
  output [15:0] io_deq_bits_1,
  output [15:0] io_deq_bits_2,
  output [15:0] io_deq_bits_3,
  output [15:0] io_deq_bits_4,
  output [15:0] io_deq_bits_5,
  output [15:0] io_deq_bits_6,
  output [15:0] io_deq_bits_7
);
  reg [15:0] _T__0 [0:3]; // @[Decoupled.scala 215:24]
  reg [31:0] _RAND_0;
  wire [15:0] _T__0__T_18_data; // @[Decoupled.scala 215:24]
  wire [1:0] _T__0__T_18_addr; // @[Decoupled.scala 215:24]
  wire [15:0] _T__0__T_10_data; // @[Decoupled.scala 215:24]
  wire [1:0] _T__0__T_10_addr; // @[Decoupled.scala 215:24]
  wire  _T__0__T_10_mask; // @[Decoupled.scala 215:24]
  wire  _T__0__T_10_en; // @[Decoupled.scala 215:24]
  reg [15:0] _T__1 [0:3]; // @[Decoupled.scala 215:24]
  reg [31:0] _RAND_1;
  wire [15:0] _T__1__T_18_data; // @[Decoupled.scala 215:24]
  wire [1:0] _T__1__T_18_addr; // @[Decoupled.scala 215:24]
  wire [15:0] _T__1__T_10_data; // @[Decoupled.scala 215:24]
  wire [1:0] _T__1__T_10_addr; // @[Decoupled.scala 215:24]
  wire  _T__1__T_10_mask; // @[Decoupled.scala 215:24]
  wire  _T__1__T_10_en; // @[Decoupled.scala 215:24]
  reg [15:0] _T__2 [0:3]; // @[Decoupled.scala 215:24]
  reg [31:0] _RAND_2;
  wire [15:0] _T__2__T_18_data; // @[Decoupled.scala 215:24]
  wire [1:0] _T__2__T_18_addr; // @[Decoupled.scala 215:24]
  wire [15:0] _T__2__T_10_data; // @[Decoupled.scala 215:24]
  wire [1:0] _T__2__T_10_addr; // @[Decoupled.scala 215:24]
  wire  _T__2__T_10_mask; // @[Decoupled.scala 215:24]
  wire  _T__2__T_10_en; // @[Decoupled.scala 215:24]
  reg [15:0] _T__3 [0:3]; // @[Decoupled.scala 215:24]
  reg [31:0] _RAND_3;
  wire [15:0] _T__3__T_18_data; // @[Decoupled.scala 215:24]
  wire [1:0] _T__3__T_18_addr; // @[Decoupled.scala 215:24]
  wire [15:0] _T__3__T_10_data; // @[Decoupled.scala 215:24]
  wire [1:0] _T__3__T_10_addr; // @[Decoupled.scala 215:24]
  wire  _T__3__T_10_mask; // @[Decoupled.scala 215:24]
  wire  _T__3__T_10_en; // @[Decoupled.scala 215:24]
  reg [15:0] _T__4 [0:3]; // @[Decoupled.scala 215:24]
  reg [31:0] _RAND_4;
  wire [15:0] _T__4__T_18_data; // @[Decoupled.scala 215:24]
  wire [1:0] _T__4__T_18_addr; // @[Decoupled.scala 215:24]
  wire [15:0] _T__4__T_10_data; // @[Decoupled.scala 215:24]
  wire [1:0] _T__4__T_10_addr; // @[Decoupled.scala 215:24]
  wire  _T__4__T_10_mask; // @[Decoupled.scala 215:24]
  wire  _T__4__T_10_en; // @[Decoupled.scala 215:24]
  reg [15:0] _T__5 [0:3]; // @[Decoupled.scala 215:24]
  reg [31:0] _RAND_5;
  wire [15:0] _T__5__T_18_data; // @[Decoupled.scala 215:24]
  wire [1:0] _T__5__T_18_addr; // @[Decoupled.scala 215:24]
  wire [15:0] _T__5__T_10_data; // @[Decoupled.scala 215:24]
  wire [1:0] _T__5__T_10_addr; // @[Decoupled.scala 215:24]
  wire  _T__5__T_10_mask; // @[Decoupled.scala 215:24]
  wire  _T__5__T_10_en; // @[Decoupled.scala 215:24]
  reg [15:0] _T__6 [0:3]; // @[Decoupled.scala 215:24]
  reg [31:0] _RAND_6;
  wire [15:0] _T__6__T_18_data; // @[Decoupled.scala 215:24]
  wire [1:0] _T__6__T_18_addr; // @[Decoupled.scala 215:24]
  wire [15:0] _T__6__T_10_data; // @[Decoupled.scala 215:24]
  wire [1:0] _T__6__T_10_addr; // @[Decoupled.scala 215:24]
  wire  _T__6__T_10_mask; // @[Decoupled.scala 215:24]
  wire  _T__6__T_10_en; // @[Decoupled.scala 215:24]
  reg [15:0] _T__7 [0:3]; // @[Decoupled.scala 215:24]
  reg [31:0] _RAND_7;
  wire [15:0] _T__7__T_18_data; // @[Decoupled.scala 215:24]
  wire [1:0] _T__7__T_18_addr; // @[Decoupled.scala 215:24]
  wire [15:0] _T__7__T_10_data; // @[Decoupled.scala 215:24]
  wire [1:0] _T__7__T_10_addr; // @[Decoupled.scala 215:24]
  wire  _T__7__T_10_mask; // @[Decoupled.scala 215:24]
  wire  _T__7__T_10_en; // @[Decoupled.scala 215:24]
  reg [1:0] value; // @[Counter.scala 26:33]
  reg [31:0] _RAND_8;
  reg [1:0] value_1; // @[Counter.scala 26:33]
  reg [31:0] _RAND_9;
  reg  _T_1; // @[Decoupled.scala 218:35]
  reg [31:0] _RAND_10;
  wire  _T_2; // @[Decoupled.scala 220:41]
  wire  _T_3; // @[Decoupled.scala 221:36]
  wire  _T_4; // @[Decoupled.scala 221:33]
  wire  _T_5; // @[Decoupled.scala 222:32]
  wire  _T_6; // @[Decoupled.scala 37:37]
  wire  _T_8; // @[Decoupled.scala 37:37]
  wire [1:0] _T_12; // @[Counter.scala 35:22]
  wire [1:0] _T_14; // @[Counter.scala 35:22]
  wire  _T_15; // @[Decoupled.scala 233:16]
  wire  _T_17; // @[Decoupled.scala 238:19]
  assign _T__0__T_18_addr = value_1;
  assign _T__0__T_18_data = _T__0[_T__0__T_18_addr]; // @[Decoupled.scala 215:24]
  assign _T__0__T_10_data = io_enq_bits_0;
  assign _T__0__T_10_addr = value;
  assign _T__0__T_10_mask = 1'h1;
  assign _T__0__T_10_en = io_enq_ready & io_enq_valid;
  assign _T__1__T_18_addr = value_1;
  assign _T__1__T_18_data = _T__1[_T__1__T_18_addr]; // @[Decoupled.scala 215:24]
  assign _T__1__T_10_data = io_enq_bits_1;
  assign _T__1__T_10_addr = value;
  assign _T__1__T_10_mask = 1'h1;
  assign _T__1__T_10_en = io_enq_ready & io_enq_valid;
  assign _T__2__T_18_addr = value_1;
  assign _T__2__T_18_data = _T__2[_T__2__T_18_addr]; // @[Decoupled.scala 215:24]
  assign _T__2__T_10_data = io_enq_bits_2;
  assign _T__2__T_10_addr = value;
  assign _T__2__T_10_mask = 1'h1;
  assign _T__2__T_10_en = io_enq_ready & io_enq_valid;
  assign _T__3__T_18_addr = value_1;
  assign _T__3__T_18_data = _T__3[_T__3__T_18_addr]; // @[Decoupled.scala 215:24]
  assign _T__3__T_10_data = io_enq_bits_3;
  assign _T__3__T_10_addr = value;
  assign _T__3__T_10_mask = 1'h1;
  assign _T__3__T_10_en = io_enq_ready & io_enq_valid;
  assign _T__4__T_18_addr = value_1;
  assign _T__4__T_18_data = _T__4[_T__4__T_18_addr]; // @[Decoupled.scala 215:24]
  assign _T__4__T_10_data = io_enq_bits_4;
  assign _T__4__T_10_addr = value;
  assign _T__4__T_10_mask = 1'h1;
  assign _T__4__T_10_en = io_enq_ready & io_enq_valid;
  assign _T__5__T_18_addr = value_1;
  assign _T__5__T_18_data = _T__5[_T__5__T_18_addr]; // @[Decoupled.scala 215:24]
  assign _T__5__T_10_data = io_enq_bits_5;
  assign _T__5__T_10_addr = value;
  assign _T__5__T_10_mask = 1'h1;
  assign _T__5__T_10_en = io_enq_ready & io_enq_valid;
  assign _T__6__T_18_addr = value_1;
  assign _T__6__T_18_data = _T__6[_T__6__T_18_addr]; // @[Decoupled.scala 215:24]
  assign _T__6__T_10_data = io_enq_bits_6;
  assign _T__6__T_10_addr = value;
  assign _T__6__T_10_mask = 1'h1;
  assign _T__6__T_10_en = io_enq_ready & io_enq_valid;
  assign _T__7__T_18_addr = value_1;
  assign _T__7__T_18_data = _T__7[_T__7__T_18_addr]; // @[Decoupled.scala 215:24]
  assign _T__7__T_10_data = io_enq_bits_7;
  assign _T__7__T_10_addr = value;
  assign _T__7__T_10_mask = 1'h1;
  assign _T__7__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_2 = value == value_1; // @[Decoupled.scala 220:41]
  assign _T_3 = _T_1 == 1'h0; // @[Decoupled.scala 221:36]
  assign _T_4 = _T_2 & _T_3; // @[Decoupled.scala 221:33]
  assign _T_5 = _T_2 & _T_1; // @[Decoupled.scala 222:32]
  assign _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 37:37]
  assign _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 37:37]
  assign _T_12 = value + 2'h1; // @[Counter.scala 35:22]
  assign _T_14 = value_1 + 2'h1; // @[Counter.scala 35:22]
  assign _T_15 = _T_6 != _T_8; // @[Decoupled.scala 233:16]
  assign _T_17 = _T_5 == 1'h0; // @[Decoupled.scala 238:19]
  assign io_enq_ready = io_deq_ready ? 1'h1 : _T_17; // @[Decoupled.scala 238:16 Decoupled.scala 251:40]
  assign io_deq_valid = _T_4 == 1'h0; // @[Decoupled.scala 237:16]
  assign io_deq_bits_0 = _T__0__T_18_data; // @[Decoupled.scala 239:15]
  assign io_deq_bits_1 = _T__1__T_18_data; // @[Decoupled.scala 239:15]
  assign io_deq_bits_2 = _T__2__T_18_data; // @[Decoupled.scala 239:15]
  assign io_deq_bits_3 = _T__3__T_18_data; // @[Decoupled.scala 239:15]
  assign io_deq_bits_4 = _T__4__T_18_data; // @[Decoupled.scala 239:15]
  assign io_deq_bits_5 = _T__5__T_18_data; // @[Decoupled.scala 239:15]
  assign io_deq_bits_6 = _T__6__T_18_data; // @[Decoupled.scala 239:15]
  assign io_deq_bits_7 = _T__7__T_18_data; // @[Decoupled.scala 239:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _T__0[initvar] = _RAND_0[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _T__1[initvar] = _RAND_1[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _T__2[initvar] = _RAND_2[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _T__3[initvar] = _RAND_3[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _T__4[initvar] = _RAND_4[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _T__5[initvar] = _RAND_5[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_6 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _T__6[initvar] = _RAND_6[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_7 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _T__7[initvar] = _RAND_7[15:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  value = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  value_1 = _RAND_9[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_1 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(_T__0__T_10_en & _T__0__T_10_mask) begin
      _T__0[_T__0__T_10_addr] <= _T__0__T_10_data; // @[Decoupled.scala 215:24]
    end
    if(_T__1__T_10_en & _T__1__T_10_mask) begin
      _T__1[_T__1__T_10_addr] <= _T__1__T_10_data; // @[Decoupled.scala 215:24]
    end
    if(_T__2__T_10_en & _T__2__T_10_mask) begin
      _T__2[_T__2__T_10_addr] <= _T__2__T_10_data; // @[Decoupled.scala 215:24]
    end
    if(_T__3__T_10_en & _T__3__T_10_mask) begin
      _T__3[_T__3__T_10_addr] <= _T__3__T_10_data; // @[Decoupled.scala 215:24]
    end
    if(_T__4__T_10_en & _T__4__T_10_mask) begin
      _T__4[_T__4__T_10_addr] <= _T__4__T_10_data; // @[Decoupled.scala 215:24]
    end
    if(_T__5__T_10_en & _T__5__T_10_mask) begin
      _T__5[_T__5__T_10_addr] <= _T__5__T_10_data; // @[Decoupled.scala 215:24]
    end
    if(_T__6__T_10_en & _T__6__T_10_mask) begin
      _T__6[_T__6__T_10_addr] <= _T__6__T_10_data; // @[Decoupled.scala 215:24]
    end
    if(_T__7__T_10_en & _T__7__T_10_mask) begin
      _T__7[_T__7__T_10_addr] <= _T__7__T_10_data; // @[Decoupled.scala 215:24]
    end
    if (reset) begin
      value <= 2'h0;
    end else begin
      if (_T_6) begin
        value <= _T_12;
      end
    end
    if (reset) begin
      value_1 <= 2'h0;
    end else begin
      if (_T_8) begin
        value_1 <= _T_14;
      end
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else begin
      if (_T_15) begin
        _T_1 <= _T_6;
      end
    end
  end
endmodule
module DecoupledStage_2(
  input         clock,
  input         reset,
  output        io_inp_ready,
  input         io_inp_valid,
  input  [15:0] io_inp_bits_0,
  input  [15:0] io_inp_bits_1,
  input  [15:0] io_inp_bits_2,
  input  [15:0] io_inp_bits_3,
  input  [15:0] io_inp_bits_4,
  input  [15:0] io_inp_bits_5,
  input  [15:0] io_inp_bits_6,
  input  [15:0] io_inp_bits_7,
  input         io_out_ready,
  output        io_out_valid,
  output [15:0] io_out_bits_0,
  output [15:0] io_out_bits_1,
  output [15:0] io_out_bits_2,
  output [15:0] io_out_bits_3,
  output [15:0] io_out_bits_4,
  output [15:0] io_out_bits_5,
  output [15:0] io_out_bits_6,
  output [15:0] io_out_bits_7
);
  reg  out_valid; // @[DecoupledStage.scala 14:22]
  reg [31:0] _RAND_0;
  reg [15:0] out_bits_0; // @[DecoupledStage.scala 15:21]
  reg [31:0] _RAND_1;
  reg [15:0] out_bits_1; // @[DecoupledStage.scala 15:21]
  reg [31:0] _RAND_2;
  reg [15:0] out_bits_2; // @[DecoupledStage.scala 15:21]
  reg [31:0] _RAND_3;
  reg [15:0] out_bits_3; // @[DecoupledStage.scala 15:21]
  reg [31:0] _RAND_4;
  reg [15:0] out_bits_4; // @[DecoupledStage.scala 15:21]
  reg [31:0] _RAND_5;
  reg [15:0] out_bits_5; // @[DecoupledStage.scala 15:21]
  reg [31:0] _RAND_6;
  reg [15:0] out_bits_6; // @[DecoupledStage.scala 15:21]
  reg [31:0] _RAND_7;
  reg [15:0] out_bits_7; // @[DecoupledStage.scala 15:21]
  reg [31:0] _RAND_8;
  wire  _T; // @[DecoupledStage.scala 20:34]
  wire  _T_2; // @[DecoupledStage.scala 22:31]
  wire  _T_3; // @[DecoupledStage.scala 22:29]
  assign _T = ~ io_out_valid; // @[DecoupledStage.scala 20:34]
  assign _T_2 = ~ io_inp_ready; // @[DecoupledStage.scala 22:31]
  assign _T_3 = io_inp_valid | _T_2; // @[DecoupledStage.scala 22:29]
  assign io_inp_ready = io_out_ready | _T; // @[DecoupledStage.scala 20:16]
  assign io_out_valid = out_valid; // @[DecoupledStage.scala 17:16]
  assign io_out_bits_0 = out_bits_0; // @[DecoupledStage.scala 18:16]
  assign io_out_bits_1 = out_bits_1; // @[DecoupledStage.scala 18:16]
  assign io_out_bits_2 = out_bits_2; // @[DecoupledStage.scala 18:16]
  assign io_out_bits_3 = out_bits_3; // @[DecoupledStage.scala 18:16]
  assign io_out_bits_4 = out_bits_4; // @[DecoupledStage.scala 18:16]
  assign io_out_bits_5 = out_bits_5; // @[DecoupledStage.scala 18:16]
  assign io_out_bits_6 = out_bits_6; // @[DecoupledStage.scala 18:16]
  assign io_out_bits_7 = out_bits_7; // @[DecoupledStage.scala 18:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  out_valid = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  out_bits_0 = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  out_bits_1 = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_bits_2 = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_bits_3 = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  out_bits_4 = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  out_bits_5 = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  out_bits_6 = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  out_bits_7 = _RAND_8[15:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      out_valid <= 1'h0;
    end else begin
      out_valid <= _T_3;
    end
    if (io_inp_ready) begin
      out_bits_0 <= io_inp_bits_0;
    end
    if (io_inp_ready) begin
      out_bits_1 <= io_inp_bits_1;
    end
    if (io_inp_ready) begin
      out_bits_2 <= io_inp_bits_2;
    end
    if (io_inp_ready) begin
      out_bits_3 <= io_inp_bits_3;
    end
    if (io_inp_ready) begin
      out_bits_4 <= io_inp_bits_4;
    end
    if (io_inp_ready) begin
      out_bits_5 <= io_inp_bits_5;
    end
    if (io_inp_ready) begin
      out_bits_6 <= io_inp_bits_6;
    end
    if (io_inp_ready) begin
      out_bits_7 <= io_inp_bits_7;
    end
  end
endmodule
module Clamper(
  input         clock,
  input         reset,
  input         io_start,
  output        io_out_ready,
  input         io_out_valid,
  input  [15:0] io_out_bits_0,
  input  [15:0] io_out_bits_1,
  input  [15:0] io_out_bits_2,
  input  [15:0] io_out_bits_3,
  input  [15:0] io_out_bits_4,
  input  [15:0] io_out_bits_5,
  input  [15:0] io_out_bits_6,
  input  [15:0] io_out_bits_7,
  input         io_res_ready,
  output        io_res_valid,
  output [15:0] io_res_bits_0,
  output [15:0] io_res_bits_1,
  output [15:0] io_res_bits_2,
  output [15:0] io_res_bits_3,
  output [15:0] io_res_bits_4,
  output [15:0] io_res_bits_5,
  output [15:0] io_res_bits_6,
  output [15:0] io_res_bits_7
);
  wire  splitOut_io_start; // @[Clamper.scala 209:24]
  wire  splitOut_io_out_ready; // @[Clamper.scala 209:24]
  wire  splitOut_io_out_valid; // @[Clamper.scala 209:24]
  wire [15:0] splitOut_io_out_bits_0; // @[Clamper.scala 209:24]
  wire [15:0] splitOut_io_out_bits_1; // @[Clamper.scala 209:24]
  wire [15:0] splitOut_io_out_bits_2; // @[Clamper.scala 209:24]
  wire [15:0] splitOut_io_out_bits_3; // @[Clamper.scala 209:24]
  wire [15:0] splitOut_io_out_bits_4; // @[Clamper.scala 209:24]
  wire [15:0] splitOut_io_out_bits_5; // @[Clamper.scala 209:24]
  wire [15:0] splitOut_io_out_bits_6; // @[Clamper.scala 209:24]
  wire [15:0] splitOut_io_out_bits_7; // @[Clamper.scala 209:24]
  wire  splitOut_io_out0_ready; // @[Clamper.scala 209:24]
  wire  splitOut_io_out0_valid; // @[Clamper.scala 209:24]
  wire [15:0] splitOut_io_out0_bits_0; // @[Clamper.scala 209:24]
  wire [15:0] splitOut_io_out0_bits_1; // @[Clamper.scala 209:24]
  wire [15:0] splitOut_io_out0_bits_2; // @[Clamper.scala 209:24]
  wire [15:0] splitOut_io_out0_bits_3; // @[Clamper.scala 209:24]
  wire [15:0] splitOut_io_out0_bits_4; // @[Clamper.scala 209:24]
  wire [15:0] splitOut_io_out0_bits_5; // @[Clamper.scala 209:24]
  wire [15:0] splitOut_io_out0_bits_6; // @[Clamper.scala 209:24]
  wire [15:0] splitOut_io_out0_bits_7; // @[Clamper.scala 209:24]
  wire  splitOut_io_out1_ready; // @[Clamper.scala 209:24]
  wire  splitOut_io_out1_valid; // @[Clamper.scala 209:24]
  wire [15:0] splitOut_io_out1_bits_0; // @[Clamper.scala 209:24]
  wire [15:0] splitOut_io_out1_bits_1; // @[Clamper.scala 209:24]
  wire [15:0] splitOut_io_out1_bits_2; // @[Clamper.scala 209:24]
  wire [15:0] splitOut_io_out1_bits_3; // @[Clamper.scala 209:24]
  wire [15:0] splitOut_io_out1_bits_4; // @[Clamper.scala 209:24]
  wire [15:0] splitOut_io_out1_bits_5; // @[Clamper.scala 209:24]
  wire [15:0] splitOut_io_out1_bits_6; // @[Clamper.scala 209:24]
  wire [15:0] splitOut_io_out1_bits_7; // @[Clamper.scala 209:24]
  wire  computeBest_clock; // @[Clamper.scala 210:27]
  wire  computeBest_reset; // @[Clamper.scala 210:27]
  wire  computeBest_io_start; // @[Clamper.scala 210:27]
  wire  computeBest_io_out0_ready; // @[Clamper.scala 210:27]
  wire  computeBest_io_out0_valid; // @[Clamper.scala 210:27]
  wire [15:0] computeBest_io_out0_bits_0; // @[Clamper.scala 210:27]
  wire [15:0] computeBest_io_out0_bits_1; // @[Clamper.scala 210:27]
  wire [15:0] computeBest_io_out0_bits_2; // @[Clamper.scala 210:27]
  wire [15:0] computeBest_io_out0_bits_3; // @[Clamper.scala 210:27]
  wire [15:0] computeBest_io_out0_bits_4; // @[Clamper.scala 210:27]
  wire [15:0] computeBest_io_out0_bits_5; // @[Clamper.scala 210:27]
  wire [15:0] computeBest_io_out0_bits_6; // @[Clamper.scala 210:27]
  wire [15:0] computeBest_io_out0_bits_7; // @[Clamper.scala 210:27]
  wire  computeBest_io_obest_ready; // @[Clamper.scala 210:27]
  wire  computeBest_io_obest_valid; // @[Clamper.scala 210:27]
  wire [15:0] computeBest_io_obest_bits; // @[Clamper.scala 210:27]
  wire  subtractOut_clock; // @[Clamper.scala 211:27]
  wire  subtractOut_reset; // @[Clamper.scala 211:27]
  wire  subtractOut_io_start; // @[Clamper.scala 211:27]
  wire  subtractOut_io_out1_ready; // @[Clamper.scala 211:27]
  wire  subtractOut_io_out1_valid; // @[Clamper.scala 211:27]
  wire [15:0] subtractOut_io_out1_bits_0; // @[Clamper.scala 211:27]
  wire [15:0] subtractOut_io_out1_bits_1; // @[Clamper.scala 211:27]
  wire [15:0] subtractOut_io_out1_bits_2; // @[Clamper.scala 211:27]
  wire [15:0] subtractOut_io_out1_bits_3; // @[Clamper.scala 211:27]
  wire [15:0] subtractOut_io_out1_bits_4; // @[Clamper.scala 211:27]
  wire [15:0] subtractOut_io_out1_bits_5; // @[Clamper.scala 211:27]
  wire [15:0] subtractOut_io_out1_bits_6; // @[Clamper.scala 211:27]
  wire [15:0] subtractOut_io_out1_bits_7; // @[Clamper.scala 211:27]
  wire  subtractOut_io_obest_ready; // @[Clamper.scala 211:27]
  wire  subtractOut_io_obest_valid; // @[Clamper.scala 211:27]
  wire [15:0] subtractOut_io_obest_bits; // @[Clamper.scala 211:27]
  wire  subtractOut_io_res_ready; // @[Clamper.scala 211:27]
  wire  subtractOut_io_res_valid; // @[Clamper.scala 211:27]
  wire [15:0] subtractOut_io_res_bits_0; // @[Clamper.scala 211:27]
  wire [15:0] subtractOut_io_res_bits_1; // @[Clamper.scala 211:27]
  wire [15:0] subtractOut_io_res_bits_2; // @[Clamper.scala 211:27]
  wire [15:0] subtractOut_io_res_bits_3; // @[Clamper.scala 211:27]
  wire [15:0] subtractOut_io_res_bits_4; // @[Clamper.scala 211:27]
  wire [15:0] subtractOut_io_res_bits_5; // @[Clamper.scala 211:27]
  wire [15:0] subtractOut_io_res_bits_6; // @[Clamper.scala 211:27]
  wire [15:0] subtractOut_io_res_bits_7; // @[Clamper.scala 211:27]
  wire  DecoupledStage_clock; // @[DecoupledStage.scala 30:19]
  wire  DecoupledStage_reset; // @[DecoupledStage.scala 30:19]
  wire  DecoupledStage_io_inp_ready; // @[DecoupledStage.scala 30:19]
  wire  DecoupledStage_io_inp_valid; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_io_inp_bits_0; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_io_inp_bits_1; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_io_inp_bits_2; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_io_inp_bits_3; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_io_inp_bits_4; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_io_inp_bits_5; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_io_inp_bits_6; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_io_inp_bits_7; // @[DecoupledStage.scala 30:19]
  wire  DecoupledStage_io_out_ready; // @[DecoupledStage.scala 30:19]
  wire  DecoupledStage_io_out_valid; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_io_out_bits_0; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_io_out_bits_1; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_io_out_bits_2; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_io_out_bits_3; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_io_out_bits_4; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_io_out_bits_5; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_io_out_bits_6; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_io_out_bits_7; // @[DecoupledStage.scala 30:19]
  wire  DecoupledStage_1_clock; // @[DecoupledStage.scala 30:19]
  wire  DecoupledStage_1_reset; // @[DecoupledStage.scala 30:19]
  wire  DecoupledStage_1_io_inp_ready; // @[DecoupledStage.scala 30:19]
  wire  DecoupledStage_1_io_inp_valid; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_1_io_inp_bits; // @[DecoupledStage.scala 30:19]
  wire  DecoupledStage_1_io_out_ready; // @[DecoupledStage.scala 30:19]
  wire  DecoupledStage_1_io_out_valid; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_1_io_out_bits; // @[DecoupledStage.scala 30:19]
  wire  Queue_clock; // @[Decoupled.scala 294:21]
  wire  Queue_reset; // @[Decoupled.scala 294:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 294:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 294:21]
  wire [15:0] Queue_io_enq_bits_0; // @[Decoupled.scala 294:21]
  wire [15:0] Queue_io_enq_bits_1; // @[Decoupled.scala 294:21]
  wire [15:0] Queue_io_enq_bits_2; // @[Decoupled.scala 294:21]
  wire [15:0] Queue_io_enq_bits_3; // @[Decoupled.scala 294:21]
  wire [15:0] Queue_io_enq_bits_4; // @[Decoupled.scala 294:21]
  wire [15:0] Queue_io_enq_bits_5; // @[Decoupled.scala 294:21]
  wire [15:0] Queue_io_enq_bits_6; // @[Decoupled.scala 294:21]
  wire [15:0] Queue_io_enq_bits_7; // @[Decoupled.scala 294:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 294:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 294:21]
  wire [15:0] Queue_io_deq_bits_0; // @[Decoupled.scala 294:21]
  wire [15:0] Queue_io_deq_bits_1; // @[Decoupled.scala 294:21]
  wire [15:0] Queue_io_deq_bits_2; // @[Decoupled.scala 294:21]
  wire [15:0] Queue_io_deq_bits_3; // @[Decoupled.scala 294:21]
  wire [15:0] Queue_io_deq_bits_4; // @[Decoupled.scala 294:21]
  wire [15:0] Queue_io_deq_bits_5; // @[Decoupled.scala 294:21]
  wire [15:0] Queue_io_deq_bits_6; // @[Decoupled.scala 294:21]
  wire [15:0] Queue_io_deq_bits_7; // @[Decoupled.scala 294:21]
  wire  DecoupledStage_2_clock; // @[DecoupledStage.scala 30:19]
  wire  DecoupledStage_2_reset; // @[DecoupledStage.scala 30:19]
  wire  DecoupledStage_2_io_inp_ready; // @[DecoupledStage.scala 30:19]
  wire  DecoupledStage_2_io_inp_valid; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_2_io_inp_bits_0; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_2_io_inp_bits_1; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_2_io_inp_bits_2; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_2_io_inp_bits_3; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_2_io_inp_bits_4; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_2_io_inp_bits_5; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_2_io_inp_bits_6; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_2_io_inp_bits_7; // @[DecoupledStage.scala 30:19]
  wire  DecoupledStage_2_io_out_ready; // @[DecoupledStage.scala 30:19]
  wire  DecoupledStage_2_io_out_valid; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_2_io_out_bits_0; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_2_io_out_bits_1; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_2_io_out_bits_2; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_2_io_out_bits_3; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_2_io_out_bits_4; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_2_io_out_bits_5; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_2_io_out_bits_6; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_2_io_out_bits_7; // @[DecoupledStage.scala 30:19]
  SplitOut splitOut ( // @[Clamper.scala 209:24]
    .io_start(splitOut_io_start),
    .io_out_ready(splitOut_io_out_ready),
    .io_out_valid(splitOut_io_out_valid),
    .io_out_bits_0(splitOut_io_out_bits_0),
    .io_out_bits_1(splitOut_io_out_bits_1),
    .io_out_bits_2(splitOut_io_out_bits_2),
    .io_out_bits_3(splitOut_io_out_bits_3),
    .io_out_bits_4(splitOut_io_out_bits_4),
    .io_out_bits_5(splitOut_io_out_bits_5),
    .io_out_bits_6(splitOut_io_out_bits_6),
    .io_out_bits_7(splitOut_io_out_bits_7),
    .io_out0_ready(splitOut_io_out0_ready),
    .io_out0_valid(splitOut_io_out0_valid),
    .io_out0_bits_0(splitOut_io_out0_bits_0),
    .io_out0_bits_1(splitOut_io_out0_bits_1),
    .io_out0_bits_2(splitOut_io_out0_bits_2),
    .io_out0_bits_3(splitOut_io_out0_bits_3),
    .io_out0_bits_4(splitOut_io_out0_bits_4),
    .io_out0_bits_5(splitOut_io_out0_bits_5),
    .io_out0_bits_6(splitOut_io_out0_bits_6),
    .io_out0_bits_7(splitOut_io_out0_bits_7),
    .io_out1_ready(splitOut_io_out1_ready),
    .io_out1_valid(splitOut_io_out1_valid),
    .io_out1_bits_0(splitOut_io_out1_bits_0),
    .io_out1_bits_1(splitOut_io_out1_bits_1),
    .io_out1_bits_2(splitOut_io_out1_bits_2),
    .io_out1_bits_3(splitOut_io_out1_bits_3),
    .io_out1_bits_4(splitOut_io_out1_bits_4),
    .io_out1_bits_5(splitOut_io_out1_bits_5),
    .io_out1_bits_6(splitOut_io_out1_bits_6),
    .io_out1_bits_7(splitOut_io_out1_bits_7)
  );
  ComputeBest computeBest ( // @[Clamper.scala 210:27]
    .clock(computeBest_clock),
    .reset(computeBest_reset),
    .io_start(computeBest_io_start),
    .io_out0_ready(computeBest_io_out0_ready),
    .io_out0_valid(computeBest_io_out0_valid),
    .io_out0_bits_0(computeBest_io_out0_bits_0),
    .io_out0_bits_1(computeBest_io_out0_bits_1),
    .io_out0_bits_2(computeBest_io_out0_bits_2),
    .io_out0_bits_3(computeBest_io_out0_bits_3),
    .io_out0_bits_4(computeBest_io_out0_bits_4),
    .io_out0_bits_5(computeBest_io_out0_bits_5),
    .io_out0_bits_6(computeBest_io_out0_bits_6),
    .io_out0_bits_7(computeBest_io_out0_bits_7),
    .io_obest_ready(computeBest_io_obest_ready),
    .io_obest_valid(computeBest_io_obest_valid),
    .io_obest_bits(computeBest_io_obest_bits)
  );
  SubtractOut subtractOut ( // @[Clamper.scala 211:27]
    .clock(subtractOut_clock),
    .reset(subtractOut_reset),
    .io_start(subtractOut_io_start),
    .io_out1_ready(subtractOut_io_out1_ready),
    .io_out1_valid(subtractOut_io_out1_valid),
    .io_out1_bits_0(subtractOut_io_out1_bits_0),
    .io_out1_bits_1(subtractOut_io_out1_bits_1),
    .io_out1_bits_2(subtractOut_io_out1_bits_2),
    .io_out1_bits_3(subtractOut_io_out1_bits_3),
    .io_out1_bits_4(subtractOut_io_out1_bits_4),
    .io_out1_bits_5(subtractOut_io_out1_bits_5),
    .io_out1_bits_6(subtractOut_io_out1_bits_6),
    .io_out1_bits_7(subtractOut_io_out1_bits_7),
    .io_obest_ready(subtractOut_io_obest_ready),
    .io_obest_valid(subtractOut_io_obest_valid),
    .io_obest_bits(subtractOut_io_obest_bits),
    .io_res_ready(subtractOut_io_res_ready),
    .io_res_valid(subtractOut_io_res_valid),
    .io_res_bits_0(subtractOut_io_res_bits_0),
    .io_res_bits_1(subtractOut_io_res_bits_1),
    .io_res_bits_2(subtractOut_io_res_bits_2),
    .io_res_bits_3(subtractOut_io_res_bits_3),
    .io_res_bits_4(subtractOut_io_res_bits_4),
    .io_res_bits_5(subtractOut_io_res_bits_5),
    .io_res_bits_6(subtractOut_io_res_bits_6),
    .io_res_bits_7(subtractOut_io_res_bits_7)
  );
  DecoupledStage DecoupledStage ( // @[DecoupledStage.scala 30:19]
    .clock(DecoupledStage_clock),
    .reset(DecoupledStage_reset),
    .io_inp_ready(DecoupledStage_io_inp_ready),
    .io_inp_valid(DecoupledStage_io_inp_valid),
    .io_inp_bits_0(DecoupledStage_io_inp_bits_0),
    .io_inp_bits_1(DecoupledStage_io_inp_bits_1),
    .io_inp_bits_2(DecoupledStage_io_inp_bits_2),
    .io_inp_bits_3(DecoupledStage_io_inp_bits_3),
    .io_inp_bits_4(DecoupledStage_io_inp_bits_4),
    .io_inp_bits_5(DecoupledStage_io_inp_bits_5),
    .io_inp_bits_6(DecoupledStage_io_inp_bits_6),
    .io_inp_bits_7(DecoupledStage_io_inp_bits_7),
    .io_out_ready(DecoupledStage_io_out_ready),
    .io_out_valid(DecoupledStage_io_out_valid),
    .io_out_bits_0(DecoupledStage_io_out_bits_0),
    .io_out_bits_1(DecoupledStage_io_out_bits_1),
    .io_out_bits_2(DecoupledStage_io_out_bits_2),
    .io_out_bits_3(DecoupledStage_io_out_bits_3),
    .io_out_bits_4(DecoupledStage_io_out_bits_4),
    .io_out_bits_5(DecoupledStage_io_out_bits_5),
    .io_out_bits_6(DecoupledStage_io_out_bits_6),
    .io_out_bits_7(DecoupledStage_io_out_bits_7)
  );
  DecoupledStage_1 DecoupledStage_1 ( // @[DecoupledStage.scala 30:19]
    .clock(DecoupledStage_1_clock),
    .reset(DecoupledStage_1_reset),
    .io_inp_ready(DecoupledStage_1_io_inp_ready),
    .io_inp_valid(DecoupledStage_1_io_inp_valid),
    .io_inp_bits(DecoupledStage_1_io_inp_bits),
    .io_out_ready(DecoupledStage_1_io_out_ready),
    .io_out_valid(DecoupledStage_1_io_out_valid),
    .io_out_bits(DecoupledStage_1_io_out_bits)
  );
  Queue Queue ( // @[Decoupled.scala 294:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_0(Queue_io_enq_bits_0),
    .io_enq_bits_1(Queue_io_enq_bits_1),
    .io_enq_bits_2(Queue_io_enq_bits_2),
    .io_enq_bits_3(Queue_io_enq_bits_3),
    .io_enq_bits_4(Queue_io_enq_bits_4),
    .io_enq_bits_5(Queue_io_enq_bits_5),
    .io_enq_bits_6(Queue_io_enq_bits_6),
    .io_enq_bits_7(Queue_io_enq_bits_7),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_0(Queue_io_deq_bits_0),
    .io_deq_bits_1(Queue_io_deq_bits_1),
    .io_deq_bits_2(Queue_io_deq_bits_2),
    .io_deq_bits_3(Queue_io_deq_bits_3),
    .io_deq_bits_4(Queue_io_deq_bits_4),
    .io_deq_bits_5(Queue_io_deq_bits_5),
    .io_deq_bits_6(Queue_io_deq_bits_6),
    .io_deq_bits_7(Queue_io_deq_bits_7)
  );
  DecoupledStage_2 DecoupledStage_2 ( // @[DecoupledStage.scala 30:19]
    .clock(DecoupledStage_2_clock),
    .reset(DecoupledStage_2_reset),
    .io_inp_ready(DecoupledStage_2_io_inp_ready),
    .io_inp_valid(DecoupledStage_2_io_inp_valid),
    .io_inp_bits_0(DecoupledStage_2_io_inp_bits_0),
    .io_inp_bits_1(DecoupledStage_2_io_inp_bits_1),
    .io_inp_bits_2(DecoupledStage_2_io_inp_bits_2),
    .io_inp_bits_3(DecoupledStage_2_io_inp_bits_3),
    .io_inp_bits_4(DecoupledStage_2_io_inp_bits_4),
    .io_inp_bits_5(DecoupledStage_2_io_inp_bits_5),
    .io_inp_bits_6(DecoupledStage_2_io_inp_bits_6),
    .io_inp_bits_7(DecoupledStage_2_io_inp_bits_7),
    .io_out_ready(DecoupledStage_2_io_out_ready),
    .io_out_valid(DecoupledStage_2_io_out_valid),
    .io_out_bits_0(DecoupledStage_2_io_out_bits_0),
    .io_out_bits_1(DecoupledStage_2_io_out_bits_1),
    .io_out_bits_2(DecoupledStage_2_io_out_bits_2),
    .io_out_bits_3(DecoupledStage_2_io_out_bits_3),
    .io_out_bits_4(DecoupledStage_2_io_out_bits_4),
    .io_out_bits_5(DecoupledStage_2_io_out_bits_5),
    .io_out_bits_6(DecoupledStage_2_io_out_bits_6),
    .io_out_bits_7(DecoupledStage_2_io_out_bits_7)
  );
  assign io_out_ready = splitOut_io_out_ready; // @[Clamper.scala 213:19]
  assign io_res_valid = DecoupledStage_2_io_out_valid; // @[Clamper.scala 223:10]
  assign io_res_bits_0 = DecoupledStage_2_io_out_bits_0; // @[Clamper.scala 223:10]
  assign io_res_bits_1 = DecoupledStage_2_io_out_bits_1; // @[Clamper.scala 223:10]
  assign io_res_bits_2 = DecoupledStage_2_io_out_bits_2; // @[Clamper.scala 223:10]
  assign io_res_bits_3 = DecoupledStage_2_io_out_bits_3; // @[Clamper.scala 223:10]
  assign io_res_bits_4 = DecoupledStage_2_io_out_bits_4; // @[Clamper.scala 223:10]
  assign io_res_bits_5 = DecoupledStage_2_io_out_bits_5; // @[Clamper.scala 223:10]
  assign io_res_bits_6 = DecoupledStage_2_io_out_bits_6; // @[Clamper.scala 223:10]
  assign io_res_bits_7 = DecoupledStage_2_io_out_bits_7; // @[Clamper.scala 223:10]
  assign splitOut_io_start = io_start; // @[Clamper.scala 214:21]
  assign splitOut_io_out_valid = io_out_valid; // @[Clamper.scala 213:19]
  assign splitOut_io_out_bits_0 = io_out_bits_0; // @[Clamper.scala 213:19]
  assign splitOut_io_out_bits_1 = io_out_bits_1; // @[Clamper.scala 213:19]
  assign splitOut_io_out_bits_2 = io_out_bits_2; // @[Clamper.scala 213:19]
  assign splitOut_io_out_bits_3 = io_out_bits_3; // @[Clamper.scala 213:19]
  assign splitOut_io_out_bits_4 = io_out_bits_4; // @[Clamper.scala 213:19]
  assign splitOut_io_out_bits_5 = io_out_bits_5; // @[Clamper.scala 213:19]
  assign splitOut_io_out_bits_6 = io_out_bits_6; // @[Clamper.scala 213:19]
  assign splitOut_io_out_bits_7 = io_out_bits_7; // @[Clamper.scala 213:19]
  assign splitOut_io_out0_ready = DecoupledStage_io_inp_ready; // @[DecoupledStage.scala 33:15]
  assign splitOut_io_out1_ready = Queue_io_enq_ready; // @[Decoupled.scala 297:17]
  assign computeBest_clock = clock;
  assign computeBest_reset = reset;
  assign computeBest_io_start = io_start; // @[Clamper.scala 217:24]
  assign computeBest_io_out0_valid = DecoupledStage_io_out_valid; // @[Clamper.scala 216:23]
  assign computeBest_io_out0_bits_0 = DecoupledStage_io_out_bits_0; // @[Clamper.scala 216:23]
  assign computeBest_io_out0_bits_1 = DecoupledStage_io_out_bits_1; // @[Clamper.scala 216:23]
  assign computeBest_io_out0_bits_2 = DecoupledStage_io_out_bits_2; // @[Clamper.scala 216:23]
  assign computeBest_io_out0_bits_3 = DecoupledStage_io_out_bits_3; // @[Clamper.scala 216:23]
  assign computeBest_io_out0_bits_4 = DecoupledStage_io_out_bits_4; // @[Clamper.scala 216:23]
  assign computeBest_io_out0_bits_5 = DecoupledStage_io_out_bits_5; // @[Clamper.scala 216:23]
  assign computeBest_io_out0_bits_6 = DecoupledStage_io_out_bits_6; // @[Clamper.scala 216:23]
  assign computeBest_io_out0_bits_7 = DecoupledStage_io_out_bits_7; // @[Clamper.scala 216:23]
  assign computeBest_io_obest_ready = DecoupledStage_1_io_inp_ready; // @[DecoupledStage.scala 33:15]
  assign subtractOut_clock = clock;
  assign subtractOut_reset = reset;
  assign subtractOut_io_start = io_start; // @[Clamper.scala 221:24]
  assign subtractOut_io_out1_valid = Queue_io_deq_valid; // @[Clamper.scala 220:23]
  assign subtractOut_io_out1_bits_0 = Queue_io_deq_bits_0; // @[Clamper.scala 220:23]
  assign subtractOut_io_out1_bits_1 = Queue_io_deq_bits_1; // @[Clamper.scala 220:23]
  assign subtractOut_io_out1_bits_2 = Queue_io_deq_bits_2; // @[Clamper.scala 220:23]
  assign subtractOut_io_out1_bits_3 = Queue_io_deq_bits_3; // @[Clamper.scala 220:23]
  assign subtractOut_io_out1_bits_4 = Queue_io_deq_bits_4; // @[Clamper.scala 220:23]
  assign subtractOut_io_out1_bits_5 = Queue_io_deq_bits_5; // @[Clamper.scala 220:23]
  assign subtractOut_io_out1_bits_6 = Queue_io_deq_bits_6; // @[Clamper.scala 220:23]
  assign subtractOut_io_out1_bits_7 = Queue_io_deq_bits_7; // @[Clamper.scala 220:23]
  assign subtractOut_io_obest_valid = DecoupledStage_1_io_out_valid; // @[Clamper.scala 219:24]
  assign subtractOut_io_obest_bits = DecoupledStage_1_io_out_bits; // @[Clamper.scala 219:24]
  assign subtractOut_io_res_ready = DecoupledStage_2_io_inp_ready; // @[DecoupledStage.scala 33:15]
  assign DecoupledStage_clock = clock;
  assign DecoupledStage_reset = reset;
  assign DecoupledStage_io_inp_valid = splitOut_io_out0_valid; // @[DecoupledStage.scala 31:20]
  assign DecoupledStage_io_inp_bits_0 = splitOut_io_out0_bits_0; // @[DecoupledStage.scala 32:19]
  assign DecoupledStage_io_inp_bits_1 = splitOut_io_out0_bits_1; // @[DecoupledStage.scala 32:19]
  assign DecoupledStage_io_inp_bits_2 = splitOut_io_out0_bits_2; // @[DecoupledStage.scala 32:19]
  assign DecoupledStage_io_inp_bits_3 = splitOut_io_out0_bits_3; // @[DecoupledStage.scala 32:19]
  assign DecoupledStage_io_inp_bits_4 = splitOut_io_out0_bits_4; // @[DecoupledStage.scala 32:19]
  assign DecoupledStage_io_inp_bits_5 = splitOut_io_out0_bits_5; // @[DecoupledStage.scala 32:19]
  assign DecoupledStage_io_inp_bits_6 = splitOut_io_out0_bits_6; // @[DecoupledStage.scala 32:19]
  assign DecoupledStage_io_inp_bits_7 = splitOut_io_out0_bits_7; // @[DecoupledStage.scala 32:19]
  assign DecoupledStage_io_out_ready = computeBest_io_out0_ready; // @[Clamper.scala 216:23]
  assign DecoupledStage_1_clock = clock;
  assign DecoupledStage_1_reset = reset;
  assign DecoupledStage_1_io_inp_valid = computeBest_io_obest_valid; // @[DecoupledStage.scala 31:20]
  assign DecoupledStage_1_io_inp_bits = computeBest_io_obest_bits; // @[DecoupledStage.scala 32:19]
  assign DecoupledStage_1_io_out_ready = subtractOut_io_obest_ready; // @[Clamper.scala 219:24]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = splitOut_io_out1_valid; // @[Decoupled.scala 295:22]
  assign Queue_io_enq_bits_0 = splitOut_io_out1_bits_0; // @[Decoupled.scala 296:21]
  assign Queue_io_enq_bits_1 = splitOut_io_out1_bits_1; // @[Decoupled.scala 296:21]
  assign Queue_io_enq_bits_2 = splitOut_io_out1_bits_2; // @[Decoupled.scala 296:21]
  assign Queue_io_enq_bits_3 = splitOut_io_out1_bits_3; // @[Decoupled.scala 296:21]
  assign Queue_io_enq_bits_4 = splitOut_io_out1_bits_4; // @[Decoupled.scala 296:21]
  assign Queue_io_enq_bits_5 = splitOut_io_out1_bits_5; // @[Decoupled.scala 296:21]
  assign Queue_io_enq_bits_6 = splitOut_io_out1_bits_6; // @[Decoupled.scala 296:21]
  assign Queue_io_enq_bits_7 = splitOut_io_out1_bits_7; // @[Decoupled.scala 296:21]
  assign Queue_io_deq_ready = subtractOut_io_out1_ready; // @[Clamper.scala 220:23]
  assign DecoupledStage_2_clock = clock;
  assign DecoupledStage_2_reset = reset;
  assign DecoupledStage_2_io_inp_valid = subtractOut_io_res_valid; // @[DecoupledStage.scala 31:20]
  assign DecoupledStage_2_io_inp_bits_0 = subtractOut_io_res_bits_0; // @[DecoupledStage.scala 32:19]
  assign DecoupledStage_2_io_inp_bits_1 = subtractOut_io_res_bits_1; // @[DecoupledStage.scala 32:19]
  assign DecoupledStage_2_io_inp_bits_2 = subtractOut_io_res_bits_2; // @[DecoupledStage.scala 32:19]
  assign DecoupledStage_2_io_inp_bits_3 = subtractOut_io_res_bits_3; // @[DecoupledStage.scala 32:19]
  assign DecoupledStage_2_io_inp_bits_4 = subtractOut_io_res_bits_4; // @[DecoupledStage.scala 32:19]
  assign DecoupledStage_2_io_inp_bits_5 = subtractOut_io_res_bits_5; // @[DecoupledStage.scala 32:19]
  assign DecoupledStage_2_io_inp_bits_6 = subtractOut_io_res_bits_6; // @[DecoupledStage.scala 32:19]
  assign DecoupledStage_2_io_inp_bits_7 = subtractOut_io_res_bits_7; // @[DecoupledStage.scala 32:19]
  assign DecoupledStage_2_io_out_ready = io_res_ready; // @[Clamper.scala 223:10]
endmodule
module Queue_1(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [15:0] io_enq_bits_0,
  input  [15:0] io_enq_bits_1,
  input  [15:0] io_enq_bits_2,
  input  [15:0] io_enq_bits_3,
  input  [15:0] io_enq_bits_4,
  input  [15:0] io_enq_bits_5,
  input  [15:0] io_enq_bits_6,
  input  [15:0] io_enq_bits_7,
  input         io_deq_ready,
  output        io_deq_valid,
  output [15:0] io_deq_bits_0,
  output [15:0] io_deq_bits_1,
  output [15:0] io_deq_bits_2,
  output [15:0] io_deq_bits_3,
  output [15:0] io_deq_bits_4,
  output [15:0] io_deq_bits_5,
  output [15:0] io_deq_bits_6,
  output [15:0] io_deq_bits_7
);
  reg [15:0] _T__0 [0:127]; // @[Decoupled.scala 215:24]
  reg [31:0] _RAND_0;
  wire [15:0] _T__0__T_18_data; // @[Decoupled.scala 215:24]
  wire [6:0] _T__0__T_18_addr; // @[Decoupled.scala 215:24]
  wire [15:0] _T__0__T_10_data; // @[Decoupled.scala 215:24]
  wire [6:0] _T__0__T_10_addr; // @[Decoupled.scala 215:24]
  wire  _T__0__T_10_mask; // @[Decoupled.scala 215:24]
  wire  _T__0__T_10_en; // @[Decoupled.scala 215:24]
  reg [15:0] _T__1 [0:127]; // @[Decoupled.scala 215:24]
  reg [31:0] _RAND_1;
  wire [15:0] _T__1__T_18_data; // @[Decoupled.scala 215:24]
  wire [6:0] _T__1__T_18_addr; // @[Decoupled.scala 215:24]
  wire [15:0] _T__1__T_10_data; // @[Decoupled.scala 215:24]
  wire [6:0] _T__1__T_10_addr; // @[Decoupled.scala 215:24]
  wire  _T__1__T_10_mask; // @[Decoupled.scala 215:24]
  wire  _T__1__T_10_en; // @[Decoupled.scala 215:24]
  reg [15:0] _T__2 [0:127]; // @[Decoupled.scala 215:24]
  reg [31:0] _RAND_2;
  wire [15:0] _T__2__T_18_data; // @[Decoupled.scala 215:24]
  wire [6:0] _T__2__T_18_addr; // @[Decoupled.scala 215:24]
  wire [15:0] _T__2__T_10_data; // @[Decoupled.scala 215:24]
  wire [6:0] _T__2__T_10_addr; // @[Decoupled.scala 215:24]
  wire  _T__2__T_10_mask; // @[Decoupled.scala 215:24]
  wire  _T__2__T_10_en; // @[Decoupled.scala 215:24]
  reg [15:0] _T__3 [0:127]; // @[Decoupled.scala 215:24]
  reg [31:0] _RAND_3;
  wire [15:0] _T__3__T_18_data; // @[Decoupled.scala 215:24]
  wire [6:0] _T__3__T_18_addr; // @[Decoupled.scala 215:24]
  wire [15:0] _T__3__T_10_data; // @[Decoupled.scala 215:24]
  wire [6:0] _T__3__T_10_addr; // @[Decoupled.scala 215:24]
  wire  _T__3__T_10_mask; // @[Decoupled.scala 215:24]
  wire  _T__3__T_10_en; // @[Decoupled.scala 215:24]
  reg [15:0] _T__4 [0:127]; // @[Decoupled.scala 215:24]
  reg [31:0] _RAND_4;
  wire [15:0] _T__4__T_18_data; // @[Decoupled.scala 215:24]
  wire [6:0] _T__4__T_18_addr; // @[Decoupled.scala 215:24]
  wire [15:0] _T__4__T_10_data; // @[Decoupled.scala 215:24]
  wire [6:0] _T__4__T_10_addr; // @[Decoupled.scala 215:24]
  wire  _T__4__T_10_mask; // @[Decoupled.scala 215:24]
  wire  _T__4__T_10_en; // @[Decoupled.scala 215:24]
  reg [15:0] _T__5 [0:127]; // @[Decoupled.scala 215:24]
  reg [31:0] _RAND_5;
  wire [15:0] _T__5__T_18_data; // @[Decoupled.scala 215:24]
  wire [6:0] _T__5__T_18_addr; // @[Decoupled.scala 215:24]
  wire [15:0] _T__5__T_10_data; // @[Decoupled.scala 215:24]
  wire [6:0] _T__5__T_10_addr; // @[Decoupled.scala 215:24]
  wire  _T__5__T_10_mask; // @[Decoupled.scala 215:24]
  wire  _T__5__T_10_en; // @[Decoupled.scala 215:24]
  reg [15:0] _T__6 [0:127]; // @[Decoupled.scala 215:24]
  reg [31:0] _RAND_6;
  wire [15:0] _T__6__T_18_data; // @[Decoupled.scala 215:24]
  wire [6:0] _T__6__T_18_addr; // @[Decoupled.scala 215:24]
  wire [15:0] _T__6__T_10_data; // @[Decoupled.scala 215:24]
  wire [6:0] _T__6__T_10_addr; // @[Decoupled.scala 215:24]
  wire  _T__6__T_10_mask; // @[Decoupled.scala 215:24]
  wire  _T__6__T_10_en; // @[Decoupled.scala 215:24]
  reg [15:0] _T__7 [0:127]; // @[Decoupled.scala 215:24]
  reg [31:0] _RAND_7;
  wire [15:0] _T__7__T_18_data; // @[Decoupled.scala 215:24]
  wire [6:0] _T__7__T_18_addr; // @[Decoupled.scala 215:24]
  wire [15:0] _T__7__T_10_data; // @[Decoupled.scala 215:24]
  wire [6:0] _T__7__T_10_addr; // @[Decoupled.scala 215:24]
  wire  _T__7__T_10_mask; // @[Decoupled.scala 215:24]
  wire  _T__7__T_10_en; // @[Decoupled.scala 215:24]
  reg [6:0] value; // @[Counter.scala 26:33]
  reg [31:0] _RAND_8;
  reg [6:0] value_1; // @[Counter.scala 26:33]
  reg [31:0] _RAND_9;
  reg  _T_1; // @[Decoupled.scala 218:35]
  reg [31:0] _RAND_10;
  wire  _T_2; // @[Decoupled.scala 220:41]
  wire  _T_3; // @[Decoupled.scala 221:36]
  wire  _T_4; // @[Decoupled.scala 221:33]
  wire  _T_5; // @[Decoupled.scala 222:32]
  wire  _T_6; // @[Decoupled.scala 37:37]
  wire  _T_8; // @[Decoupled.scala 37:37]
  wire [6:0] _T_12; // @[Counter.scala 35:22]
  wire [6:0] _T_14; // @[Counter.scala 35:22]
  wire  _T_15; // @[Decoupled.scala 233:16]
  wire  _T_17; // @[Decoupled.scala 238:19]
  assign _T__0__T_18_addr = value_1;
  assign _T__0__T_18_data = _T__0[_T__0__T_18_addr]; // @[Decoupled.scala 215:24]
  assign _T__0__T_10_data = io_enq_bits_0;
  assign _T__0__T_10_addr = value;
  assign _T__0__T_10_mask = 1'h1;
  assign _T__0__T_10_en = io_enq_ready & io_enq_valid;
  assign _T__1__T_18_addr = value_1;
  assign _T__1__T_18_data = _T__1[_T__1__T_18_addr]; // @[Decoupled.scala 215:24]
  assign _T__1__T_10_data = io_enq_bits_1;
  assign _T__1__T_10_addr = value;
  assign _T__1__T_10_mask = 1'h1;
  assign _T__1__T_10_en = io_enq_ready & io_enq_valid;
  assign _T__2__T_18_addr = value_1;
  assign _T__2__T_18_data = _T__2[_T__2__T_18_addr]; // @[Decoupled.scala 215:24]
  assign _T__2__T_10_data = io_enq_bits_2;
  assign _T__2__T_10_addr = value;
  assign _T__2__T_10_mask = 1'h1;
  assign _T__2__T_10_en = io_enq_ready & io_enq_valid;
  assign _T__3__T_18_addr = value_1;
  assign _T__3__T_18_data = _T__3[_T__3__T_18_addr]; // @[Decoupled.scala 215:24]
  assign _T__3__T_10_data = io_enq_bits_3;
  assign _T__3__T_10_addr = value;
  assign _T__3__T_10_mask = 1'h1;
  assign _T__3__T_10_en = io_enq_ready & io_enq_valid;
  assign _T__4__T_18_addr = value_1;
  assign _T__4__T_18_data = _T__4[_T__4__T_18_addr]; // @[Decoupled.scala 215:24]
  assign _T__4__T_10_data = io_enq_bits_4;
  assign _T__4__T_10_addr = value;
  assign _T__4__T_10_mask = 1'h1;
  assign _T__4__T_10_en = io_enq_ready & io_enq_valid;
  assign _T__5__T_18_addr = value_1;
  assign _T__5__T_18_data = _T__5[_T__5__T_18_addr]; // @[Decoupled.scala 215:24]
  assign _T__5__T_10_data = io_enq_bits_5;
  assign _T__5__T_10_addr = value;
  assign _T__5__T_10_mask = 1'h1;
  assign _T__5__T_10_en = io_enq_ready & io_enq_valid;
  assign _T__6__T_18_addr = value_1;
  assign _T__6__T_18_data = _T__6[_T__6__T_18_addr]; // @[Decoupled.scala 215:24]
  assign _T__6__T_10_data = io_enq_bits_6;
  assign _T__6__T_10_addr = value;
  assign _T__6__T_10_mask = 1'h1;
  assign _T__6__T_10_en = io_enq_ready & io_enq_valid;
  assign _T__7__T_18_addr = value_1;
  assign _T__7__T_18_data = _T__7[_T__7__T_18_addr]; // @[Decoupled.scala 215:24]
  assign _T__7__T_10_data = io_enq_bits_7;
  assign _T__7__T_10_addr = value;
  assign _T__7__T_10_mask = 1'h1;
  assign _T__7__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_2 = value == value_1; // @[Decoupled.scala 220:41]
  assign _T_3 = _T_1 == 1'h0; // @[Decoupled.scala 221:36]
  assign _T_4 = _T_2 & _T_3; // @[Decoupled.scala 221:33]
  assign _T_5 = _T_2 & _T_1; // @[Decoupled.scala 222:32]
  assign _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 37:37]
  assign _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 37:37]
  assign _T_12 = value + 7'h1; // @[Counter.scala 35:22]
  assign _T_14 = value_1 + 7'h1; // @[Counter.scala 35:22]
  assign _T_15 = _T_6 != _T_8; // @[Decoupled.scala 233:16]
  assign _T_17 = _T_5 == 1'h0; // @[Decoupled.scala 238:19]
  assign io_enq_ready = io_deq_ready ? 1'h1 : _T_17; // @[Decoupled.scala 238:16 Decoupled.scala 251:40]
  assign io_deq_valid = _T_4 == 1'h0; // @[Decoupled.scala 237:16]
  assign io_deq_bits_0 = _T__0__T_18_data; // @[Decoupled.scala 239:15]
  assign io_deq_bits_1 = _T__1__T_18_data; // @[Decoupled.scala 239:15]
  assign io_deq_bits_2 = _T__2__T_18_data; // @[Decoupled.scala 239:15]
  assign io_deq_bits_3 = _T__3__T_18_data; // @[Decoupled.scala 239:15]
  assign io_deq_bits_4 = _T__4__T_18_data; // @[Decoupled.scala 239:15]
  assign io_deq_bits_5 = _T__5__T_18_data; // @[Decoupled.scala 239:15]
  assign io_deq_bits_6 = _T__6__T_18_data; // @[Decoupled.scala 239:15]
  assign io_deq_bits_7 = _T__7__T_18_data; // @[Decoupled.scala 239:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    _T__0[initvar] = _RAND_0[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    _T__1[initvar] = _RAND_1[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    _T__2[initvar] = _RAND_2[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    _T__3[initvar] = _RAND_3[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    _T__4[initvar] = _RAND_4[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    _T__5[initvar] = _RAND_5[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_6 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    _T__6[initvar] = _RAND_6[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_7 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    _T__7[initvar] = _RAND_7[15:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  value = _RAND_8[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  value_1 = _RAND_9[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_1 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(_T__0__T_10_en & _T__0__T_10_mask) begin
      _T__0[_T__0__T_10_addr] <= _T__0__T_10_data; // @[Decoupled.scala 215:24]
    end
    if(_T__1__T_10_en & _T__1__T_10_mask) begin
      _T__1[_T__1__T_10_addr] <= _T__1__T_10_data; // @[Decoupled.scala 215:24]
    end
    if(_T__2__T_10_en & _T__2__T_10_mask) begin
      _T__2[_T__2__T_10_addr] <= _T__2__T_10_data; // @[Decoupled.scala 215:24]
    end
    if(_T__3__T_10_en & _T__3__T_10_mask) begin
      _T__3[_T__3__T_10_addr] <= _T__3__T_10_data; // @[Decoupled.scala 215:24]
    end
    if(_T__4__T_10_en & _T__4__T_10_mask) begin
      _T__4[_T__4__T_10_addr] <= _T__4__T_10_data; // @[Decoupled.scala 215:24]
    end
    if(_T__5__T_10_en & _T__5__T_10_mask) begin
      _T__5[_T__5__T_10_addr] <= _T__5__T_10_data; // @[Decoupled.scala 215:24]
    end
    if(_T__6__T_10_en & _T__6__T_10_mask) begin
      _T__6[_T__6__T_10_addr] <= _T__6__T_10_data; // @[Decoupled.scala 215:24]
    end
    if(_T__7__T_10_en & _T__7__T_10_mask) begin
      _T__7[_T__7__T_10_addr] <= _T__7__T_10_data; // @[Decoupled.scala 215:24]
    end
    if (reset) begin
      value <= 7'h0;
    end else begin
      if (_T_6) begin
        value <= _T_12;
      end
    end
    if (reset) begin
      value_1 <= 7'h0;
    end else begin
      if (_T_8) begin
        value_1 <= _T_14;
      end
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else begin
      if (_T_15) begin
        _T_1 <= _T_6;
      end
    end
  end
endmodule
module Queue_2(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [15:0] io_enq_bits_0,
  input  [15:0] io_enq_bits_1,
  input  [15:0] io_enq_bits_2,
  input  [15:0] io_enq_bits_3,
  input  [15:0] io_enq_bits_4,
  input  [15:0] io_enq_bits_5,
  input  [15:0] io_enq_bits_6,
  input  [15:0] io_enq_bits_7,
  input         io_deq_ready,
  output        io_deq_valid,
  output [15:0] io_deq_bits_0,
  output [15:0] io_deq_bits_1,
  output [15:0] io_deq_bits_2,
  output [15:0] io_deq_bits_3,
  output [15:0] io_deq_bits_4,
  output [15:0] io_deq_bits_5,
  output [15:0] io_deq_bits_6,
  output [15:0] io_deq_bits_7
);
  reg [15:0] _T__0 [0:3]; // @[Decoupled.scala 215:24]
  reg [31:0] _RAND_0;
  wire [15:0] _T__0__T_18_data; // @[Decoupled.scala 215:24]
  wire [1:0] _T__0__T_18_addr; // @[Decoupled.scala 215:24]
  wire [15:0] _T__0__T_10_data; // @[Decoupled.scala 215:24]
  wire [1:0] _T__0__T_10_addr; // @[Decoupled.scala 215:24]
  wire  _T__0__T_10_mask; // @[Decoupled.scala 215:24]
  wire  _T__0__T_10_en; // @[Decoupled.scala 215:24]
  reg [15:0] _T__1 [0:3]; // @[Decoupled.scala 215:24]
  reg [31:0] _RAND_1;
  wire [15:0] _T__1__T_18_data; // @[Decoupled.scala 215:24]
  wire [1:0] _T__1__T_18_addr; // @[Decoupled.scala 215:24]
  wire [15:0] _T__1__T_10_data; // @[Decoupled.scala 215:24]
  wire [1:0] _T__1__T_10_addr; // @[Decoupled.scala 215:24]
  wire  _T__1__T_10_mask; // @[Decoupled.scala 215:24]
  wire  _T__1__T_10_en; // @[Decoupled.scala 215:24]
  reg [15:0] _T__2 [0:3]; // @[Decoupled.scala 215:24]
  reg [31:0] _RAND_2;
  wire [15:0] _T__2__T_18_data; // @[Decoupled.scala 215:24]
  wire [1:0] _T__2__T_18_addr; // @[Decoupled.scala 215:24]
  wire [15:0] _T__2__T_10_data; // @[Decoupled.scala 215:24]
  wire [1:0] _T__2__T_10_addr; // @[Decoupled.scala 215:24]
  wire  _T__2__T_10_mask; // @[Decoupled.scala 215:24]
  wire  _T__2__T_10_en; // @[Decoupled.scala 215:24]
  reg [15:0] _T__3 [0:3]; // @[Decoupled.scala 215:24]
  reg [31:0] _RAND_3;
  wire [15:0] _T__3__T_18_data; // @[Decoupled.scala 215:24]
  wire [1:0] _T__3__T_18_addr; // @[Decoupled.scala 215:24]
  wire [15:0] _T__3__T_10_data; // @[Decoupled.scala 215:24]
  wire [1:0] _T__3__T_10_addr; // @[Decoupled.scala 215:24]
  wire  _T__3__T_10_mask; // @[Decoupled.scala 215:24]
  wire  _T__3__T_10_en; // @[Decoupled.scala 215:24]
  reg [15:0] _T__4 [0:3]; // @[Decoupled.scala 215:24]
  reg [31:0] _RAND_4;
  wire [15:0] _T__4__T_18_data; // @[Decoupled.scala 215:24]
  wire [1:0] _T__4__T_18_addr; // @[Decoupled.scala 215:24]
  wire [15:0] _T__4__T_10_data; // @[Decoupled.scala 215:24]
  wire [1:0] _T__4__T_10_addr; // @[Decoupled.scala 215:24]
  wire  _T__4__T_10_mask; // @[Decoupled.scala 215:24]
  wire  _T__4__T_10_en; // @[Decoupled.scala 215:24]
  reg [15:0] _T__5 [0:3]; // @[Decoupled.scala 215:24]
  reg [31:0] _RAND_5;
  wire [15:0] _T__5__T_18_data; // @[Decoupled.scala 215:24]
  wire [1:0] _T__5__T_18_addr; // @[Decoupled.scala 215:24]
  wire [15:0] _T__5__T_10_data; // @[Decoupled.scala 215:24]
  wire [1:0] _T__5__T_10_addr; // @[Decoupled.scala 215:24]
  wire  _T__5__T_10_mask; // @[Decoupled.scala 215:24]
  wire  _T__5__T_10_en; // @[Decoupled.scala 215:24]
  reg [15:0] _T__6 [0:3]; // @[Decoupled.scala 215:24]
  reg [31:0] _RAND_6;
  wire [15:0] _T__6__T_18_data; // @[Decoupled.scala 215:24]
  wire [1:0] _T__6__T_18_addr; // @[Decoupled.scala 215:24]
  wire [15:0] _T__6__T_10_data; // @[Decoupled.scala 215:24]
  wire [1:0] _T__6__T_10_addr; // @[Decoupled.scala 215:24]
  wire  _T__6__T_10_mask; // @[Decoupled.scala 215:24]
  wire  _T__6__T_10_en; // @[Decoupled.scala 215:24]
  reg [15:0] _T__7 [0:3]; // @[Decoupled.scala 215:24]
  reg [31:0] _RAND_7;
  wire [15:0] _T__7__T_18_data; // @[Decoupled.scala 215:24]
  wire [1:0] _T__7__T_18_addr; // @[Decoupled.scala 215:24]
  wire [15:0] _T__7__T_10_data; // @[Decoupled.scala 215:24]
  wire [1:0] _T__7__T_10_addr; // @[Decoupled.scala 215:24]
  wire  _T__7__T_10_mask; // @[Decoupled.scala 215:24]
  wire  _T__7__T_10_en; // @[Decoupled.scala 215:24]
  reg [1:0] value; // @[Counter.scala 26:33]
  reg [31:0] _RAND_8;
  reg [1:0] value_1; // @[Counter.scala 26:33]
  reg [31:0] _RAND_9;
  reg  _T_1; // @[Decoupled.scala 218:35]
  reg [31:0] _RAND_10;
  wire  _T_2; // @[Decoupled.scala 220:41]
  wire  _T_3; // @[Decoupled.scala 221:36]
  wire  _T_4; // @[Decoupled.scala 221:33]
  wire  _T_5; // @[Decoupled.scala 222:32]
  wire  _T_6; // @[Decoupled.scala 37:37]
  wire  _T_8; // @[Decoupled.scala 37:37]
  wire [1:0] _T_12; // @[Counter.scala 35:22]
  wire [1:0] _T_14; // @[Counter.scala 35:22]
  wire  _T_15; // @[Decoupled.scala 233:16]
  assign _T__0__T_18_addr = value_1;
  assign _T__0__T_18_data = _T__0[_T__0__T_18_addr]; // @[Decoupled.scala 215:24]
  assign _T__0__T_10_data = io_enq_bits_0;
  assign _T__0__T_10_addr = value;
  assign _T__0__T_10_mask = 1'h1;
  assign _T__0__T_10_en = io_enq_ready & io_enq_valid;
  assign _T__1__T_18_addr = value_1;
  assign _T__1__T_18_data = _T__1[_T__1__T_18_addr]; // @[Decoupled.scala 215:24]
  assign _T__1__T_10_data = io_enq_bits_1;
  assign _T__1__T_10_addr = value;
  assign _T__1__T_10_mask = 1'h1;
  assign _T__1__T_10_en = io_enq_ready & io_enq_valid;
  assign _T__2__T_18_addr = value_1;
  assign _T__2__T_18_data = _T__2[_T__2__T_18_addr]; // @[Decoupled.scala 215:24]
  assign _T__2__T_10_data = io_enq_bits_2;
  assign _T__2__T_10_addr = value;
  assign _T__2__T_10_mask = 1'h1;
  assign _T__2__T_10_en = io_enq_ready & io_enq_valid;
  assign _T__3__T_18_addr = value_1;
  assign _T__3__T_18_data = _T__3[_T__3__T_18_addr]; // @[Decoupled.scala 215:24]
  assign _T__3__T_10_data = io_enq_bits_3;
  assign _T__3__T_10_addr = value;
  assign _T__3__T_10_mask = 1'h1;
  assign _T__3__T_10_en = io_enq_ready & io_enq_valid;
  assign _T__4__T_18_addr = value_1;
  assign _T__4__T_18_data = _T__4[_T__4__T_18_addr]; // @[Decoupled.scala 215:24]
  assign _T__4__T_10_data = io_enq_bits_4;
  assign _T__4__T_10_addr = value;
  assign _T__4__T_10_mask = 1'h1;
  assign _T__4__T_10_en = io_enq_ready & io_enq_valid;
  assign _T__5__T_18_addr = value_1;
  assign _T__5__T_18_data = _T__5[_T__5__T_18_addr]; // @[Decoupled.scala 215:24]
  assign _T__5__T_10_data = io_enq_bits_5;
  assign _T__5__T_10_addr = value;
  assign _T__5__T_10_mask = 1'h1;
  assign _T__5__T_10_en = io_enq_ready & io_enq_valid;
  assign _T__6__T_18_addr = value_1;
  assign _T__6__T_18_data = _T__6[_T__6__T_18_addr]; // @[Decoupled.scala 215:24]
  assign _T__6__T_10_data = io_enq_bits_6;
  assign _T__6__T_10_addr = value;
  assign _T__6__T_10_mask = 1'h1;
  assign _T__6__T_10_en = io_enq_ready & io_enq_valid;
  assign _T__7__T_18_addr = value_1;
  assign _T__7__T_18_data = _T__7[_T__7__T_18_addr]; // @[Decoupled.scala 215:24]
  assign _T__7__T_10_data = io_enq_bits_7;
  assign _T__7__T_10_addr = value;
  assign _T__7__T_10_mask = 1'h1;
  assign _T__7__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_2 = value == value_1; // @[Decoupled.scala 220:41]
  assign _T_3 = _T_1 == 1'h0; // @[Decoupled.scala 221:36]
  assign _T_4 = _T_2 & _T_3; // @[Decoupled.scala 221:33]
  assign _T_5 = _T_2 & _T_1; // @[Decoupled.scala 222:32]
  assign _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 37:37]
  assign _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 37:37]
  assign _T_12 = value + 2'h1; // @[Counter.scala 35:22]
  assign _T_14 = value_1 + 2'h1; // @[Counter.scala 35:22]
  assign _T_15 = _T_6 != _T_8; // @[Decoupled.scala 233:16]
  assign io_enq_ready = _T_5 == 1'h0; // @[Decoupled.scala 238:16]
  assign io_deq_valid = _T_4 == 1'h0; // @[Decoupled.scala 237:16]
  assign io_deq_bits_0 = _T__0__T_18_data; // @[Decoupled.scala 239:15]
  assign io_deq_bits_1 = _T__1__T_18_data; // @[Decoupled.scala 239:15]
  assign io_deq_bits_2 = _T__2__T_18_data; // @[Decoupled.scala 239:15]
  assign io_deq_bits_3 = _T__3__T_18_data; // @[Decoupled.scala 239:15]
  assign io_deq_bits_4 = _T__4__T_18_data; // @[Decoupled.scala 239:15]
  assign io_deq_bits_5 = _T__5__T_18_data; // @[Decoupled.scala 239:15]
  assign io_deq_bits_6 = _T__6__T_18_data; // @[Decoupled.scala 239:15]
  assign io_deq_bits_7 = _T__7__T_18_data; // @[Decoupled.scala 239:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _T__0[initvar] = _RAND_0[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _T__1[initvar] = _RAND_1[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _T__2[initvar] = _RAND_2[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _T__3[initvar] = _RAND_3[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _T__4[initvar] = _RAND_4[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _T__5[initvar] = _RAND_5[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_6 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _T__6[initvar] = _RAND_6[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_7 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _T__7[initvar] = _RAND_7[15:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  value = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  value_1 = _RAND_9[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_1 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(_T__0__T_10_en & _T__0__T_10_mask) begin
      _T__0[_T__0__T_10_addr] <= _T__0__T_10_data; // @[Decoupled.scala 215:24]
    end
    if(_T__1__T_10_en & _T__1__T_10_mask) begin
      _T__1[_T__1__T_10_addr] <= _T__1__T_10_data; // @[Decoupled.scala 215:24]
    end
    if(_T__2__T_10_en & _T__2__T_10_mask) begin
      _T__2[_T__2__T_10_addr] <= _T__2__T_10_data; // @[Decoupled.scala 215:24]
    end
    if(_T__3__T_10_en & _T__3__T_10_mask) begin
      _T__3[_T__3__T_10_addr] <= _T__3__T_10_data; // @[Decoupled.scala 215:24]
    end
    if(_T__4__T_10_en & _T__4__T_10_mask) begin
      _T__4[_T__4__T_10_addr] <= _T__4__T_10_data; // @[Decoupled.scala 215:24]
    end
    if(_T__5__T_10_en & _T__5__T_10_mask) begin
      _T__5[_T__5__T_10_addr] <= _T__5__T_10_data; // @[Decoupled.scala 215:24]
    end
    if(_T__6__T_10_en & _T__6__T_10_mask) begin
      _T__6[_T__6__T_10_addr] <= _T__6__T_10_data; // @[Decoupled.scala 215:24]
    end
    if(_T__7__T_10_en & _T__7__T_10_mask) begin
      _T__7[_T__7__T_10_addr] <= _T__7__T_10_data; // @[Decoupled.scala 215:24]
    end
    if (reset) begin
      value <= 2'h0;
    end else begin
      if (_T_6) begin
        value <= _T_12;
      end
    end
    if (reset) begin
      value_1 <= 2'h0;
    end else begin
      if (_T_8) begin
        value_1 <= _T_14;
      end
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else begin
      if (_T_15) begin
        _T_1 <= _T_6;
      end
    end
  end
endmodule
module trws(
  input         clock,
  input         reset,
  input         io_start,
  output        io_done,
  input         io_modeLoad,
  input         io_modeCompute,
  input         io_loadIdx,
  input         io_computeIdx,
  output        io_gi_ready,
  input         io_gi_valid,
  input  [15:0] io_gi_bits_0,
  input  [15:0] io_gi_bits_1,
  input  [15:0] io_gi_bits_2,
  input  [15:0] io_gi_bits_3,
  input  [15:0] io_gi_bits_4,
  input  [15:0] io_gi_bits_5,
  input  [15:0] io_gi_bits_6,
  input  [15:0] io_gi_bits_7,
  output        io_wi_ready,
  input         io_wi_valid,
  input  [15:0] io_wi_bits_0,
  input  [15:0] io_wi_bits_1,
  input  [15:0] io_wi_bits_2,
  input  [15:0] io_wi_bits_3,
  input  [15:0] io_wi_bits_4,
  input  [15:0] io_wi_bits_5,
  input  [15:0] io_wi_bits_6,
  input  [15:0] io_wi_bits_7,
  output        io_mi_ready,
  input         io_mi_valid,
  input  [15:0] io_mi_bits_0,
  input  [15:0] io_mi_bits_1,
  input  [15:0] io_mi_bits_2,
  input  [15:0] io_mi_bits_3,
  input  [15:0] io_mi_bits_4,
  input  [15:0] io_mi_bits_5,
  input  [15:0] io_mi_bits_6,
  input  [15:0] io_mi_bits_7,
  output        io_slc_ready,
  input         io_slc_valid,
  input  [15:0] io_slc_bits_e,
  input  [15:0] io_slc_bits_a,
  output        io_lof_ready,
  input         io_lof_valid,
  input  [15:0] io_lof_bits_e,
  input  [15:0] io_lof_bits_a,
  input         io_mo_ready,
  output        io_mo_valid,
  output [15:0] io_mo_bits_bits_0,
  output [15:0] io_mo_bits_bits_1,
  output [15:0] io_mo_bits_bits_2,
  output [15:0] io_mo_bits_bits_3,
  output [15:0] io_mo_bits_bits_4,
  output [15:0] io_mo_bits_bits_5,
  output [15:0] io_mo_bits_bits_6,
  output [15:0] io_mo_bits_bits_7
);
  wire  splitter_io_mi_ready; // @[trws.scala 30:24]
  wire  splitter_io_mi_valid; // @[trws.scala 30:24]
  wire [15:0] splitter_io_mi_bits_0; // @[trws.scala 30:24]
  wire [15:0] splitter_io_mi_bits_1; // @[trws.scala 30:24]
  wire [15:0] splitter_io_mi_bits_2; // @[trws.scala 30:24]
  wire [15:0] splitter_io_mi_bits_3; // @[trws.scala 30:24]
  wire [15:0] splitter_io_mi_bits_4; // @[trws.scala 30:24]
  wire [15:0] splitter_io_mi_bits_5; // @[trws.scala 30:24]
  wire [15:0] splitter_io_mi_bits_6; // @[trws.scala 30:24]
  wire [15:0] splitter_io_mi_bits_7; // @[trws.scala 30:24]
  wire  splitter_io_mi0_ready; // @[trws.scala 30:24]
  wire  splitter_io_mi0_valid; // @[trws.scala 30:24]
  wire [15:0] splitter_io_mi0_bits_0; // @[trws.scala 30:24]
  wire [15:0] splitter_io_mi0_bits_1; // @[trws.scala 30:24]
  wire [15:0] splitter_io_mi0_bits_2; // @[trws.scala 30:24]
  wire [15:0] splitter_io_mi0_bits_3; // @[trws.scala 30:24]
  wire [15:0] splitter_io_mi0_bits_4; // @[trws.scala 30:24]
  wire [15:0] splitter_io_mi0_bits_5; // @[trws.scala 30:24]
  wire [15:0] splitter_io_mi0_bits_6; // @[trws.scala 30:24]
  wire [15:0] splitter_io_mi0_bits_7; // @[trws.scala 30:24]
  wire  splitter_io_mi1_ready; // @[trws.scala 30:24]
  wire  splitter_io_mi1_valid; // @[trws.scala 30:24]
  wire [15:0] splitter_io_mi1_bits_0; // @[trws.scala 30:24]
  wire [15:0] splitter_io_mi1_bits_1; // @[trws.scala 30:24]
  wire [15:0] splitter_io_mi1_bits_2; // @[trws.scala 30:24]
  wire [15:0] splitter_io_mi1_bits_3; // @[trws.scala 30:24]
  wire [15:0] splitter_io_mi1_bits_4; // @[trws.scala 30:24]
  wire [15:0] splitter_io_mi1_bits_5; // @[trws.scala 30:24]
  wire [15:0] splitter_io_mi1_bits_6; // @[trws.scala 30:24]
  wire [15:0] splitter_io_mi1_bits_7; // @[trws.scala 30:24]
  wire  frontend_clock; // @[trws.scala 31:24]
  wire  frontend_reset; // @[trws.scala 31:24]
  wire  frontend_io_start; // @[trws.scala 31:24]
  wire  frontend_io_gi_ready; // @[trws.scala 31:24]
  wire  frontend_io_gi_valid; // @[trws.scala 31:24]
  wire [15:0] frontend_io_gi_bits_0; // @[trws.scala 31:24]
  wire [15:0] frontend_io_gi_bits_1; // @[trws.scala 31:24]
  wire [15:0] frontend_io_gi_bits_2; // @[trws.scala 31:24]
  wire [15:0] frontend_io_gi_bits_3; // @[trws.scala 31:24]
  wire [15:0] frontend_io_gi_bits_4; // @[trws.scala 31:24]
  wire [15:0] frontend_io_gi_bits_5; // @[trws.scala 31:24]
  wire [15:0] frontend_io_gi_bits_6; // @[trws.scala 31:24]
  wire [15:0] frontend_io_gi_bits_7; // @[trws.scala 31:24]
  wire  frontend_io_wi_ready; // @[trws.scala 31:24]
  wire  frontend_io_wi_valid; // @[trws.scala 31:24]
  wire [15:0] frontend_io_wi_bits_0; // @[trws.scala 31:24]
  wire [15:0] frontend_io_wi_bits_1; // @[trws.scala 31:24]
  wire [15:0] frontend_io_wi_bits_2; // @[trws.scala 31:24]
  wire [15:0] frontend_io_wi_bits_3; // @[trws.scala 31:24]
  wire [15:0] frontend_io_wi_bits_4; // @[trws.scala 31:24]
  wire [15:0] frontend_io_wi_bits_5; // @[trws.scala 31:24]
  wire [15:0] frontend_io_wi_bits_6; // @[trws.scala 31:24]
  wire [15:0] frontend_io_wi_bits_7; // @[trws.scala 31:24]
  wire  frontend_io_a0_ready; // @[trws.scala 31:24]
  wire  frontend_io_a0_valid; // @[trws.scala 31:24]
  wire [15:0] frontend_io_a0_bits_0; // @[trws.scala 31:24]
  wire [15:0] frontend_io_a0_bits_1; // @[trws.scala 31:24]
  wire [15:0] frontend_io_a0_bits_2; // @[trws.scala 31:24]
  wire [15:0] frontend_io_a0_bits_3; // @[trws.scala 31:24]
  wire [15:0] frontend_io_a0_bits_4; // @[trws.scala 31:24]
  wire [15:0] frontend_io_a0_bits_5; // @[trws.scala 31:24]
  wire [15:0] frontend_io_a0_bits_6; // @[trws.scala 31:24]
  wire [15:0] frontend_io_a0_bits_7; // @[trws.scala 31:24]
  wire  frontend_io_mi1_ready; // @[trws.scala 31:24]
  wire  frontend_io_mi1_valid; // @[trws.scala 31:24]
  wire [15:0] frontend_io_mi1_bits_0; // @[trws.scala 31:24]
  wire [15:0] frontend_io_mi1_bits_1; // @[trws.scala 31:24]
  wire [15:0] frontend_io_mi1_bits_2; // @[trws.scala 31:24]
  wire [15:0] frontend_io_mi1_bits_3; // @[trws.scala 31:24]
  wire [15:0] frontend_io_mi1_bits_4; // @[trws.scala 31:24]
  wire [15:0] frontend_io_mi1_bits_5; // @[trws.scala 31:24]
  wire [15:0] frontend_io_mi1_bits_6; // @[trws.scala 31:24]
  wire [15:0] frontend_io_mi1_bits_7; // @[trws.scala 31:24]
  wire  frontend_io_adj_ready; // @[trws.scala 31:24]
  wire  frontend_io_adj_valid; // @[trws.scala 31:24]
  wire [15:0] frontend_io_adj_bits_0; // @[trws.scala 31:24]
  wire [15:0] frontend_io_adj_bits_1; // @[trws.scala 31:24]
  wire [15:0] frontend_io_adj_bits_2; // @[trws.scala 31:24]
  wire [15:0] frontend_io_adj_bits_3; // @[trws.scala 31:24]
  wire [15:0] frontend_io_adj_bits_4; // @[trws.scala 31:24]
  wire [15:0] frontend_io_adj_bits_5; // @[trws.scala 31:24]
  wire [15:0] frontend_io_adj_bits_6; // @[trws.scala 31:24]
  wire [15:0] frontend_io_adj_bits_7; // @[trws.scala 31:24]
  wire  frontend_io_off_ready; // @[trws.scala 31:24]
  wire  frontend_io_off_valid; // @[trws.scala 31:24]
  wire [15:0] frontend_io_off_bits_0; // @[trws.scala 31:24]
  wire [15:0] frontend_io_off_bits_1; // @[trws.scala 31:24]
  wire [15:0] frontend_io_off_bits_2; // @[trws.scala 31:24]
  wire [15:0] frontend_io_off_bits_3; // @[trws.scala 31:24]
  wire [15:0] frontend_io_off_bits_4; // @[trws.scala 31:24]
  wire [15:0] frontend_io_off_bits_5; // @[trws.scala 31:24]
  wire [15:0] frontend_io_off_bits_6; // @[trws.scala 31:24]
  wire [15:0] frontend_io_off_bits_7; // @[trws.scala 31:24]
  wire  backend_clock; // @[trws.scala 32:23]
  wire  backend_reset; // @[trws.scala 32:23]
  wire  backend_io_start; // @[trws.scala 32:23]
  wire  backend_io_done; // @[trws.scala 32:23]
  wire  backend_io_res_ready; // @[trws.scala 32:23]
  wire  backend_io_res_valid; // @[trws.scala 32:23]
  wire [15:0] backend_io_res_bits_0; // @[trws.scala 32:23]
  wire [15:0] backend_io_res_bits_1; // @[trws.scala 32:23]
  wire [15:0] backend_io_res_bits_2; // @[trws.scala 32:23]
  wire [15:0] backend_io_res_bits_3; // @[trws.scala 32:23]
  wire [15:0] backend_io_res_bits_4; // @[trws.scala 32:23]
  wire [15:0] backend_io_res_bits_5; // @[trws.scala 32:23]
  wire [15:0] backend_io_res_bits_6; // @[trws.scala 32:23]
  wire [15:0] backend_io_res_bits_7; // @[trws.scala 32:23]
  wire  backend_io_mo_ready; // @[trws.scala 32:23]
  wire  backend_io_mo_valid; // @[trws.scala 32:23]
  wire [15:0] backend_io_mo_bits_bits_0; // @[trws.scala 32:23]
  wire [15:0] backend_io_mo_bits_bits_1; // @[trws.scala 32:23]
  wire [15:0] backend_io_mo_bits_bits_2; // @[trws.scala 32:23]
  wire [15:0] backend_io_mo_bits_bits_3; // @[trws.scala 32:23]
  wire [15:0] backend_io_mo_bits_bits_4; // @[trws.scala 32:23]
  wire [15:0] backend_io_mo_bits_bits_5; // @[trws.scala 32:23]
  wire [15:0] backend_io_mo_bits_bits_6; // @[trws.scala 32:23]
  wire [15:0] backend_io_mo_bits_bits_7; // @[trws.scala 32:23]
  wire  backend_io_adj_ready; // @[trws.scala 32:23]
  wire  backend_io_adj_valid; // @[trws.scala 32:23]
  wire [15:0] backend_io_adj_bits_0; // @[trws.scala 32:23]
  wire [15:0] backend_io_adj_bits_1; // @[trws.scala 32:23]
  wire [15:0] backend_io_adj_bits_2; // @[trws.scala 32:23]
  wire [15:0] backend_io_adj_bits_3; // @[trws.scala 32:23]
  wire [15:0] backend_io_adj_bits_4; // @[trws.scala 32:23]
  wire [15:0] backend_io_adj_bits_5; // @[trws.scala 32:23]
  wire [15:0] backend_io_adj_bits_6; // @[trws.scala 32:23]
  wire [15:0] backend_io_adj_bits_7; // @[trws.scala 32:23]
  wire  accumulator_clock; // @[trws.scala 33:27]
  wire  accumulator_reset; // @[trws.scala 33:27]
  wire  accumulator_io_mi0_ready; // @[trws.scala 33:27]
  wire  accumulator_io_mi0_valid; // @[trws.scala 33:27]
  wire [15:0] accumulator_io_mi0_bits_0; // @[trws.scala 33:27]
  wire [15:0] accumulator_io_mi0_bits_1; // @[trws.scala 33:27]
  wire [15:0] accumulator_io_mi0_bits_2; // @[trws.scala 33:27]
  wire [15:0] accumulator_io_mi0_bits_3; // @[trws.scala 33:27]
  wire [15:0] accumulator_io_mi0_bits_4; // @[trws.scala 33:27]
  wire [15:0] accumulator_io_mi0_bits_5; // @[trws.scala 33:27]
  wire [15:0] accumulator_io_mi0_bits_6; // @[trws.scala 33:27]
  wire [15:0] accumulator_io_mi0_bits_7; // @[trws.scala 33:27]
  wire  accumulator_io_a0_ready; // @[trws.scala 33:27]
  wire  accumulator_io_a0_valid; // @[trws.scala 33:27]
  wire [15:0] accumulator_io_a0_bits_0; // @[trws.scala 33:27]
  wire [15:0] accumulator_io_a0_bits_1; // @[trws.scala 33:27]
  wire [15:0] accumulator_io_a0_bits_2; // @[trws.scala 33:27]
  wire [15:0] accumulator_io_a0_bits_3; // @[trws.scala 33:27]
  wire [15:0] accumulator_io_a0_bits_4; // @[trws.scala 33:27]
  wire [15:0] accumulator_io_a0_bits_5; // @[trws.scala 33:27]
  wire [15:0] accumulator_io_a0_bits_6; // @[trws.scala 33:27]
  wire [15:0] accumulator_io_a0_bits_7; // @[trws.scala 33:27]
  wire  loaf_clock; // @[trws.scala 35:20]
  wire  loaf_reset; // @[trws.scala 35:20]
  wire  loaf_io_start; // @[trws.scala 35:20]
  wire  loaf_io_doneLoading; // @[trws.scala 35:20]
  wire  loaf_io_modeLoad; // @[trws.scala 35:20]
  wire  loaf_io_modeCompute; // @[trws.scala 35:20]
  wire  loaf_io_loadIdx; // @[trws.scala 35:20]
  wire  loaf_io_computeIdx; // @[trws.scala 35:20]
  wire  loaf_io_off_ready; // @[trws.scala 35:20]
  wire  loaf_io_off_valid; // @[trws.scala 35:20]
  wire [15:0] loaf_io_off_bits_0; // @[trws.scala 35:20]
  wire [15:0] loaf_io_off_bits_1; // @[trws.scala 35:20]
  wire [15:0] loaf_io_off_bits_2; // @[trws.scala 35:20]
  wire [15:0] loaf_io_off_bits_3; // @[trws.scala 35:20]
  wire [15:0] loaf_io_off_bits_4; // @[trws.scala 35:20]
  wire [15:0] loaf_io_off_bits_5; // @[trws.scala 35:20]
  wire [15:0] loaf_io_off_bits_6; // @[trws.scala 35:20]
  wire [15:0] loaf_io_off_bits_7; // @[trws.scala 35:20]
  wire  loaf_io_out_ready; // @[trws.scala 35:20]
  wire  loaf_io_out_valid; // @[trws.scala 35:20]
  wire [15:0] loaf_io_out_bits_0; // @[trws.scala 35:20]
  wire [15:0] loaf_io_out_bits_1; // @[trws.scala 35:20]
  wire [15:0] loaf_io_out_bits_2; // @[trws.scala 35:20]
  wire [15:0] loaf_io_out_bits_3; // @[trws.scala 35:20]
  wire [15:0] loaf_io_out_bits_4; // @[trws.scala 35:20]
  wire [15:0] loaf_io_out_bits_5; // @[trws.scala 35:20]
  wire [15:0] loaf_io_out_bits_6; // @[trws.scala 35:20]
  wire [15:0] loaf_io_out_bits_7; // @[trws.scala 35:20]
  wire  loaf_io_slc_ready; // @[trws.scala 35:20]
  wire  loaf_io_slc_valid; // @[trws.scala 35:20]
  wire [15:0] loaf_io_slc_bits_e; // @[trws.scala 35:20]
  wire [15:0] loaf_io_slc_bits_a; // @[trws.scala 35:20]
  wire  loaf_io_lof_ready; // @[trws.scala 35:20]
  wire  loaf_io_lof_valid; // @[trws.scala 35:20]
  wire [15:0] loaf_io_lof_bits_e; // @[trws.scala 35:20]
  wire [15:0] loaf_io_lof_bits_a; // @[trws.scala 35:20]
  wire  clamper_clock; // @[trws.scala 36:23]
  wire  clamper_reset; // @[trws.scala 36:23]
  wire  clamper_io_start; // @[trws.scala 36:23]
  wire  clamper_io_out_ready; // @[trws.scala 36:23]
  wire  clamper_io_out_valid; // @[trws.scala 36:23]
  wire [15:0] clamper_io_out_bits_0; // @[trws.scala 36:23]
  wire [15:0] clamper_io_out_bits_1; // @[trws.scala 36:23]
  wire [15:0] clamper_io_out_bits_2; // @[trws.scala 36:23]
  wire [15:0] clamper_io_out_bits_3; // @[trws.scala 36:23]
  wire [15:0] clamper_io_out_bits_4; // @[trws.scala 36:23]
  wire [15:0] clamper_io_out_bits_5; // @[trws.scala 36:23]
  wire [15:0] clamper_io_out_bits_6; // @[trws.scala 36:23]
  wire [15:0] clamper_io_out_bits_7; // @[trws.scala 36:23]
  wire  clamper_io_res_ready; // @[trws.scala 36:23]
  wire  clamper_io_res_valid; // @[trws.scala 36:23]
  wire [15:0] clamper_io_res_bits_0; // @[trws.scala 36:23]
  wire [15:0] clamper_io_res_bits_1; // @[trws.scala 36:23]
  wire [15:0] clamper_io_res_bits_2; // @[trws.scala 36:23]
  wire [15:0] clamper_io_res_bits_3; // @[trws.scala 36:23]
  wire [15:0] clamper_io_res_bits_4; // @[trws.scala 36:23]
  wire [15:0] clamper_io_res_bits_5; // @[trws.scala 36:23]
  wire [15:0] clamper_io_res_bits_6; // @[trws.scala 36:23]
  wire [15:0] clamper_io_res_bits_7; // @[trws.scala 36:23]
  wire  DecoupledStage_clock; // @[DecoupledStage.scala 30:19]
  wire  DecoupledStage_reset; // @[DecoupledStage.scala 30:19]
  wire  DecoupledStage_io_inp_ready; // @[DecoupledStage.scala 30:19]
  wire  DecoupledStage_io_inp_valid; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_io_inp_bits_0; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_io_inp_bits_1; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_io_inp_bits_2; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_io_inp_bits_3; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_io_inp_bits_4; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_io_inp_bits_5; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_io_inp_bits_6; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_io_inp_bits_7; // @[DecoupledStage.scala 30:19]
  wire  DecoupledStage_io_out_ready; // @[DecoupledStage.scala 30:19]
  wire  DecoupledStage_io_out_valid; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_io_out_bits_0; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_io_out_bits_1; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_io_out_bits_2; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_io_out_bits_3; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_io_out_bits_4; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_io_out_bits_5; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_io_out_bits_6; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_io_out_bits_7; // @[DecoupledStage.scala 30:19]
  wire  DecoupledStage_1_clock; // @[DecoupledStage.scala 30:19]
  wire  DecoupledStage_1_reset; // @[DecoupledStage.scala 30:19]
  wire  DecoupledStage_1_io_inp_ready; // @[DecoupledStage.scala 30:19]
  wire  DecoupledStage_1_io_inp_valid; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_1_io_inp_bits_0; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_1_io_inp_bits_1; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_1_io_inp_bits_2; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_1_io_inp_bits_3; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_1_io_inp_bits_4; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_1_io_inp_bits_5; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_1_io_inp_bits_6; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_1_io_inp_bits_7; // @[DecoupledStage.scala 30:19]
  wire  DecoupledStage_1_io_out_ready; // @[DecoupledStage.scala 30:19]
  wire  DecoupledStage_1_io_out_valid; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_1_io_out_bits_0; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_1_io_out_bits_1; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_1_io_out_bits_2; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_1_io_out_bits_3; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_1_io_out_bits_4; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_1_io_out_bits_5; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_1_io_out_bits_6; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_1_io_out_bits_7; // @[DecoupledStage.scala 30:19]
  wire  Queue_clock; // @[Decoupled.scala 294:21]
  wire  Queue_reset; // @[Decoupled.scala 294:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 294:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 294:21]
  wire [15:0] Queue_io_enq_bits_0; // @[Decoupled.scala 294:21]
  wire [15:0] Queue_io_enq_bits_1; // @[Decoupled.scala 294:21]
  wire [15:0] Queue_io_enq_bits_2; // @[Decoupled.scala 294:21]
  wire [15:0] Queue_io_enq_bits_3; // @[Decoupled.scala 294:21]
  wire [15:0] Queue_io_enq_bits_4; // @[Decoupled.scala 294:21]
  wire [15:0] Queue_io_enq_bits_5; // @[Decoupled.scala 294:21]
  wire [15:0] Queue_io_enq_bits_6; // @[Decoupled.scala 294:21]
  wire [15:0] Queue_io_enq_bits_7; // @[Decoupled.scala 294:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 294:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 294:21]
  wire [15:0] Queue_io_deq_bits_0; // @[Decoupled.scala 294:21]
  wire [15:0] Queue_io_deq_bits_1; // @[Decoupled.scala 294:21]
  wire [15:0] Queue_io_deq_bits_2; // @[Decoupled.scala 294:21]
  wire [15:0] Queue_io_deq_bits_3; // @[Decoupled.scala 294:21]
  wire [15:0] Queue_io_deq_bits_4; // @[Decoupled.scala 294:21]
  wire [15:0] Queue_io_deq_bits_5; // @[Decoupled.scala 294:21]
  wire [15:0] Queue_io_deq_bits_6; // @[Decoupled.scala 294:21]
  wire [15:0] Queue_io_deq_bits_7; // @[Decoupled.scala 294:21]
  wire  Queue_1_clock; // @[Decoupled.scala 294:21]
  wire  Queue_1_reset; // @[Decoupled.scala 294:21]
  wire  Queue_1_io_enq_ready; // @[Decoupled.scala 294:21]
  wire  Queue_1_io_enq_valid; // @[Decoupled.scala 294:21]
  wire [15:0] Queue_1_io_enq_bits_0; // @[Decoupled.scala 294:21]
  wire [15:0] Queue_1_io_enq_bits_1; // @[Decoupled.scala 294:21]
  wire [15:0] Queue_1_io_enq_bits_2; // @[Decoupled.scala 294:21]
  wire [15:0] Queue_1_io_enq_bits_3; // @[Decoupled.scala 294:21]
  wire [15:0] Queue_1_io_enq_bits_4; // @[Decoupled.scala 294:21]
  wire [15:0] Queue_1_io_enq_bits_5; // @[Decoupled.scala 294:21]
  wire [15:0] Queue_1_io_enq_bits_6; // @[Decoupled.scala 294:21]
  wire [15:0] Queue_1_io_enq_bits_7; // @[Decoupled.scala 294:21]
  wire  Queue_1_io_deq_ready; // @[Decoupled.scala 294:21]
  wire  Queue_1_io_deq_valid; // @[Decoupled.scala 294:21]
  wire [15:0] Queue_1_io_deq_bits_0; // @[Decoupled.scala 294:21]
  wire [15:0] Queue_1_io_deq_bits_1; // @[Decoupled.scala 294:21]
  wire [15:0] Queue_1_io_deq_bits_2; // @[Decoupled.scala 294:21]
  wire [15:0] Queue_1_io_deq_bits_3; // @[Decoupled.scala 294:21]
  wire [15:0] Queue_1_io_deq_bits_4; // @[Decoupled.scala 294:21]
  wire [15:0] Queue_1_io_deq_bits_5; // @[Decoupled.scala 294:21]
  wire [15:0] Queue_1_io_deq_bits_6; // @[Decoupled.scala 294:21]
  wire [15:0] Queue_1_io_deq_bits_7; // @[Decoupled.scala 294:21]
  wire  DecoupledStage_2_clock; // @[DecoupledStage.scala 30:19]
  wire  DecoupledStage_2_reset; // @[DecoupledStage.scala 30:19]
  wire  DecoupledStage_2_io_inp_ready; // @[DecoupledStage.scala 30:19]
  wire  DecoupledStage_2_io_inp_valid; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_2_io_inp_bits_0; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_2_io_inp_bits_1; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_2_io_inp_bits_2; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_2_io_inp_bits_3; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_2_io_inp_bits_4; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_2_io_inp_bits_5; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_2_io_inp_bits_6; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_2_io_inp_bits_7; // @[DecoupledStage.scala 30:19]
  wire  DecoupledStage_2_io_out_ready; // @[DecoupledStage.scala 30:19]
  wire  DecoupledStage_2_io_out_valid; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_2_io_out_bits_0; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_2_io_out_bits_1; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_2_io_out_bits_2; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_2_io_out_bits_3; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_2_io_out_bits_4; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_2_io_out_bits_5; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_2_io_out_bits_6; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_2_io_out_bits_7; // @[DecoupledStage.scala 30:19]
  wire  DecoupledStage_3_clock; // @[DecoupledStage.scala 30:19]
  wire  DecoupledStage_3_reset; // @[DecoupledStage.scala 30:19]
  wire  DecoupledStage_3_io_inp_ready; // @[DecoupledStage.scala 30:19]
  wire  DecoupledStage_3_io_inp_valid; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_3_io_inp_bits_0; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_3_io_inp_bits_1; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_3_io_inp_bits_2; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_3_io_inp_bits_3; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_3_io_inp_bits_4; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_3_io_inp_bits_5; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_3_io_inp_bits_6; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_3_io_inp_bits_7; // @[DecoupledStage.scala 30:19]
  wire  DecoupledStage_3_io_out_ready; // @[DecoupledStage.scala 30:19]
  wire  DecoupledStage_3_io_out_valid; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_3_io_out_bits_0; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_3_io_out_bits_1; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_3_io_out_bits_2; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_3_io_out_bits_3; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_3_io_out_bits_4; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_3_io_out_bits_5; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_3_io_out_bits_6; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_3_io_out_bits_7; // @[DecoupledStage.scala 30:19]
  wire  DecoupledStage_4_clock; // @[DecoupledStage.scala 30:19]
  wire  DecoupledStage_4_reset; // @[DecoupledStage.scala 30:19]
  wire  DecoupledStage_4_io_inp_ready; // @[DecoupledStage.scala 30:19]
  wire  DecoupledStage_4_io_inp_valid; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_4_io_inp_bits_0; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_4_io_inp_bits_1; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_4_io_inp_bits_2; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_4_io_inp_bits_3; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_4_io_inp_bits_4; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_4_io_inp_bits_5; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_4_io_inp_bits_6; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_4_io_inp_bits_7; // @[DecoupledStage.scala 30:19]
  wire  DecoupledStage_4_io_out_ready; // @[DecoupledStage.scala 30:19]
  wire  DecoupledStage_4_io_out_valid; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_4_io_out_bits_0; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_4_io_out_bits_1; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_4_io_out_bits_2; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_4_io_out_bits_3; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_4_io_out_bits_4; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_4_io_out_bits_5; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_4_io_out_bits_6; // @[DecoupledStage.scala 30:19]
  wire [15:0] DecoupledStage_4_io_out_bits_7; // @[DecoupledStage.scala 30:19]
  wire  _T; // @[trws.scala 68:16]
  wire  _T_1; // @[trws.scala 68:32]
  wire  _T_2; // @[trws.scala 68:57]
  wire  _T_3; // @[trws.scala 68:70]
  Splitter splitter ( // @[trws.scala 30:24]
    .io_mi_ready(splitter_io_mi_ready),
    .io_mi_valid(splitter_io_mi_valid),
    .io_mi_bits_0(splitter_io_mi_bits_0),
    .io_mi_bits_1(splitter_io_mi_bits_1),
    .io_mi_bits_2(splitter_io_mi_bits_2),
    .io_mi_bits_3(splitter_io_mi_bits_3),
    .io_mi_bits_4(splitter_io_mi_bits_4),
    .io_mi_bits_5(splitter_io_mi_bits_5),
    .io_mi_bits_6(splitter_io_mi_bits_6),
    .io_mi_bits_7(splitter_io_mi_bits_7),
    .io_mi0_ready(splitter_io_mi0_ready),
    .io_mi0_valid(splitter_io_mi0_valid),
    .io_mi0_bits_0(splitter_io_mi0_bits_0),
    .io_mi0_bits_1(splitter_io_mi0_bits_1),
    .io_mi0_bits_2(splitter_io_mi0_bits_2),
    .io_mi0_bits_3(splitter_io_mi0_bits_3),
    .io_mi0_bits_4(splitter_io_mi0_bits_4),
    .io_mi0_bits_5(splitter_io_mi0_bits_5),
    .io_mi0_bits_6(splitter_io_mi0_bits_6),
    .io_mi0_bits_7(splitter_io_mi0_bits_7),
    .io_mi1_ready(splitter_io_mi1_ready),
    .io_mi1_valid(splitter_io_mi1_valid),
    .io_mi1_bits_0(splitter_io_mi1_bits_0),
    .io_mi1_bits_1(splitter_io_mi1_bits_1),
    .io_mi1_bits_2(splitter_io_mi1_bits_2),
    .io_mi1_bits_3(splitter_io_mi1_bits_3),
    .io_mi1_bits_4(splitter_io_mi1_bits_4),
    .io_mi1_bits_5(splitter_io_mi1_bits_5),
    .io_mi1_bits_6(splitter_io_mi1_bits_6),
    .io_mi1_bits_7(splitter_io_mi1_bits_7)
  );
  Frontend frontend ( // @[trws.scala 31:24]
    .clock(frontend_clock),
    .reset(frontend_reset),
    .io_start(frontend_io_start),
    .io_gi_ready(frontend_io_gi_ready),
    .io_gi_valid(frontend_io_gi_valid),
    .io_gi_bits_0(frontend_io_gi_bits_0),
    .io_gi_bits_1(frontend_io_gi_bits_1),
    .io_gi_bits_2(frontend_io_gi_bits_2),
    .io_gi_bits_3(frontend_io_gi_bits_3),
    .io_gi_bits_4(frontend_io_gi_bits_4),
    .io_gi_bits_5(frontend_io_gi_bits_5),
    .io_gi_bits_6(frontend_io_gi_bits_6),
    .io_gi_bits_7(frontend_io_gi_bits_7),
    .io_wi_ready(frontend_io_wi_ready),
    .io_wi_valid(frontend_io_wi_valid),
    .io_wi_bits_0(frontend_io_wi_bits_0),
    .io_wi_bits_1(frontend_io_wi_bits_1),
    .io_wi_bits_2(frontend_io_wi_bits_2),
    .io_wi_bits_3(frontend_io_wi_bits_3),
    .io_wi_bits_4(frontend_io_wi_bits_4),
    .io_wi_bits_5(frontend_io_wi_bits_5),
    .io_wi_bits_6(frontend_io_wi_bits_6),
    .io_wi_bits_7(frontend_io_wi_bits_7),
    .io_a0_ready(frontend_io_a0_ready),
    .io_a0_valid(frontend_io_a0_valid),
    .io_a0_bits_0(frontend_io_a0_bits_0),
    .io_a0_bits_1(frontend_io_a0_bits_1),
    .io_a0_bits_2(frontend_io_a0_bits_2),
    .io_a0_bits_3(frontend_io_a0_bits_3),
    .io_a0_bits_4(frontend_io_a0_bits_4),
    .io_a0_bits_5(frontend_io_a0_bits_5),
    .io_a0_bits_6(frontend_io_a0_bits_6),
    .io_a0_bits_7(frontend_io_a0_bits_7),
    .io_mi1_ready(frontend_io_mi1_ready),
    .io_mi1_valid(frontend_io_mi1_valid),
    .io_mi1_bits_0(frontend_io_mi1_bits_0),
    .io_mi1_bits_1(frontend_io_mi1_bits_1),
    .io_mi1_bits_2(frontend_io_mi1_bits_2),
    .io_mi1_bits_3(frontend_io_mi1_bits_3),
    .io_mi1_bits_4(frontend_io_mi1_bits_4),
    .io_mi1_bits_5(frontend_io_mi1_bits_5),
    .io_mi1_bits_6(frontend_io_mi1_bits_6),
    .io_mi1_bits_7(frontend_io_mi1_bits_7),
    .io_adj_ready(frontend_io_adj_ready),
    .io_adj_valid(frontend_io_adj_valid),
    .io_adj_bits_0(frontend_io_adj_bits_0),
    .io_adj_bits_1(frontend_io_adj_bits_1),
    .io_adj_bits_2(frontend_io_adj_bits_2),
    .io_adj_bits_3(frontend_io_adj_bits_3),
    .io_adj_bits_4(frontend_io_adj_bits_4),
    .io_adj_bits_5(frontend_io_adj_bits_5),
    .io_adj_bits_6(frontend_io_adj_bits_6),
    .io_adj_bits_7(frontend_io_adj_bits_7),
    .io_off_ready(frontend_io_off_ready),
    .io_off_valid(frontend_io_off_valid),
    .io_off_bits_0(frontend_io_off_bits_0),
    .io_off_bits_1(frontend_io_off_bits_1),
    .io_off_bits_2(frontend_io_off_bits_2),
    .io_off_bits_3(frontend_io_off_bits_3),
    .io_off_bits_4(frontend_io_off_bits_4),
    .io_off_bits_5(frontend_io_off_bits_5),
    .io_off_bits_6(frontend_io_off_bits_6),
    .io_off_bits_7(frontend_io_off_bits_7)
  );
  Backend backend ( // @[trws.scala 32:23]
    .clock(backend_clock),
    .reset(backend_reset),
    .io_start(backend_io_start),
    .io_done(backend_io_done),
    .io_res_ready(backend_io_res_ready),
    .io_res_valid(backend_io_res_valid),
    .io_res_bits_0(backend_io_res_bits_0),
    .io_res_bits_1(backend_io_res_bits_1),
    .io_res_bits_2(backend_io_res_bits_2),
    .io_res_bits_3(backend_io_res_bits_3),
    .io_res_bits_4(backend_io_res_bits_4),
    .io_res_bits_5(backend_io_res_bits_5),
    .io_res_bits_6(backend_io_res_bits_6),
    .io_res_bits_7(backend_io_res_bits_7),
    .io_mo_ready(backend_io_mo_ready),
    .io_mo_valid(backend_io_mo_valid),
    .io_mo_bits_bits_0(backend_io_mo_bits_bits_0),
    .io_mo_bits_bits_1(backend_io_mo_bits_bits_1),
    .io_mo_bits_bits_2(backend_io_mo_bits_bits_2),
    .io_mo_bits_bits_3(backend_io_mo_bits_bits_3),
    .io_mo_bits_bits_4(backend_io_mo_bits_bits_4),
    .io_mo_bits_bits_5(backend_io_mo_bits_bits_5),
    .io_mo_bits_bits_6(backend_io_mo_bits_bits_6),
    .io_mo_bits_bits_7(backend_io_mo_bits_bits_7),
    .io_adj_ready(backend_io_adj_ready),
    .io_adj_valid(backend_io_adj_valid),
    .io_adj_bits_0(backend_io_adj_bits_0),
    .io_adj_bits_1(backend_io_adj_bits_1),
    .io_adj_bits_2(backend_io_adj_bits_2),
    .io_adj_bits_3(backend_io_adj_bits_3),
    .io_adj_bits_4(backend_io_adj_bits_4),
    .io_adj_bits_5(backend_io_adj_bits_5),
    .io_adj_bits_6(backend_io_adj_bits_6),
    .io_adj_bits_7(backend_io_adj_bits_7)
  );
  Accumulator accumulator ( // @[trws.scala 33:27]
    .clock(accumulator_clock),
    .reset(accumulator_reset),
    .io_mi0_ready(accumulator_io_mi0_ready),
    .io_mi0_valid(accumulator_io_mi0_valid),
    .io_mi0_bits_0(accumulator_io_mi0_bits_0),
    .io_mi0_bits_1(accumulator_io_mi0_bits_1),
    .io_mi0_bits_2(accumulator_io_mi0_bits_2),
    .io_mi0_bits_3(accumulator_io_mi0_bits_3),
    .io_mi0_bits_4(accumulator_io_mi0_bits_4),
    .io_mi0_bits_5(accumulator_io_mi0_bits_5),
    .io_mi0_bits_6(accumulator_io_mi0_bits_6),
    .io_mi0_bits_7(accumulator_io_mi0_bits_7),
    .io_a0_ready(accumulator_io_a0_ready),
    .io_a0_valid(accumulator_io_a0_valid),
    .io_a0_bits_0(accumulator_io_a0_bits_0),
    .io_a0_bits_1(accumulator_io_a0_bits_1),
    .io_a0_bits_2(accumulator_io_a0_bits_2),
    .io_a0_bits_3(accumulator_io_a0_bits_3),
    .io_a0_bits_4(accumulator_io_a0_bits_4),
    .io_a0_bits_5(accumulator_io_a0_bits_5),
    .io_a0_bits_6(accumulator_io_a0_bits_6),
    .io_a0_bits_7(accumulator_io_a0_bits_7)
  );
  Loaf loaf ( // @[trws.scala 35:20]
    .clock(loaf_clock),
    .reset(loaf_reset),
    .io_start(loaf_io_start),
    .io_doneLoading(loaf_io_doneLoading),
    .io_modeLoad(loaf_io_modeLoad),
    .io_modeCompute(loaf_io_modeCompute),
    .io_loadIdx(loaf_io_loadIdx),
    .io_computeIdx(loaf_io_computeIdx),
    .io_off_ready(loaf_io_off_ready),
    .io_off_valid(loaf_io_off_valid),
    .io_off_bits_0(loaf_io_off_bits_0),
    .io_off_bits_1(loaf_io_off_bits_1),
    .io_off_bits_2(loaf_io_off_bits_2),
    .io_off_bits_3(loaf_io_off_bits_3),
    .io_off_bits_4(loaf_io_off_bits_4),
    .io_off_bits_5(loaf_io_off_bits_5),
    .io_off_bits_6(loaf_io_off_bits_6),
    .io_off_bits_7(loaf_io_off_bits_7),
    .io_out_ready(loaf_io_out_ready),
    .io_out_valid(loaf_io_out_valid),
    .io_out_bits_0(loaf_io_out_bits_0),
    .io_out_bits_1(loaf_io_out_bits_1),
    .io_out_bits_2(loaf_io_out_bits_2),
    .io_out_bits_3(loaf_io_out_bits_3),
    .io_out_bits_4(loaf_io_out_bits_4),
    .io_out_bits_5(loaf_io_out_bits_5),
    .io_out_bits_6(loaf_io_out_bits_6),
    .io_out_bits_7(loaf_io_out_bits_7),
    .io_slc_ready(loaf_io_slc_ready),
    .io_slc_valid(loaf_io_slc_valid),
    .io_slc_bits_e(loaf_io_slc_bits_e),
    .io_slc_bits_a(loaf_io_slc_bits_a),
    .io_lof_ready(loaf_io_lof_ready),
    .io_lof_valid(loaf_io_lof_valid),
    .io_lof_bits_e(loaf_io_lof_bits_e),
    .io_lof_bits_a(loaf_io_lof_bits_a)
  );
  Clamper clamper ( // @[trws.scala 36:23]
    .clock(clamper_clock),
    .reset(clamper_reset),
    .io_start(clamper_io_start),
    .io_out_ready(clamper_io_out_ready),
    .io_out_valid(clamper_io_out_valid),
    .io_out_bits_0(clamper_io_out_bits_0),
    .io_out_bits_1(clamper_io_out_bits_1),
    .io_out_bits_2(clamper_io_out_bits_2),
    .io_out_bits_3(clamper_io_out_bits_3),
    .io_out_bits_4(clamper_io_out_bits_4),
    .io_out_bits_5(clamper_io_out_bits_5),
    .io_out_bits_6(clamper_io_out_bits_6),
    .io_out_bits_7(clamper_io_out_bits_7),
    .io_res_ready(clamper_io_res_ready),
    .io_res_valid(clamper_io_res_valid),
    .io_res_bits_0(clamper_io_res_bits_0),
    .io_res_bits_1(clamper_io_res_bits_1),
    .io_res_bits_2(clamper_io_res_bits_2),
    .io_res_bits_3(clamper_io_res_bits_3),
    .io_res_bits_4(clamper_io_res_bits_4),
    .io_res_bits_5(clamper_io_res_bits_5),
    .io_res_bits_6(clamper_io_res_bits_6),
    .io_res_bits_7(clamper_io_res_bits_7)
  );
  DecoupledStage_2 DecoupledStage ( // @[DecoupledStage.scala 30:19]
    .clock(DecoupledStage_clock),
    .reset(DecoupledStage_reset),
    .io_inp_ready(DecoupledStage_io_inp_ready),
    .io_inp_valid(DecoupledStage_io_inp_valid),
    .io_inp_bits_0(DecoupledStage_io_inp_bits_0),
    .io_inp_bits_1(DecoupledStage_io_inp_bits_1),
    .io_inp_bits_2(DecoupledStage_io_inp_bits_2),
    .io_inp_bits_3(DecoupledStage_io_inp_bits_3),
    .io_inp_bits_4(DecoupledStage_io_inp_bits_4),
    .io_inp_bits_5(DecoupledStage_io_inp_bits_5),
    .io_inp_bits_6(DecoupledStage_io_inp_bits_6),
    .io_inp_bits_7(DecoupledStage_io_inp_bits_7),
    .io_out_ready(DecoupledStage_io_out_ready),
    .io_out_valid(DecoupledStage_io_out_valid),
    .io_out_bits_0(DecoupledStage_io_out_bits_0),
    .io_out_bits_1(DecoupledStage_io_out_bits_1),
    .io_out_bits_2(DecoupledStage_io_out_bits_2),
    .io_out_bits_3(DecoupledStage_io_out_bits_3),
    .io_out_bits_4(DecoupledStage_io_out_bits_4),
    .io_out_bits_5(DecoupledStage_io_out_bits_5),
    .io_out_bits_6(DecoupledStage_io_out_bits_6),
    .io_out_bits_7(DecoupledStage_io_out_bits_7)
  );
  DecoupledStage_2 DecoupledStage_1 ( // @[DecoupledStage.scala 30:19]
    .clock(DecoupledStage_1_clock),
    .reset(DecoupledStage_1_reset),
    .io_inp_ready(DecoupledStage_1_io_inp_ready),
    .io_inp_valid(DecoupledStage_1_io_inp_valid),
    .io_inp_bits_0(DecoupledStage_1_io_inp_bits_0),
    .io_inp_bits_1(DecoupledStage_1_io_inp_bits_1),
    .io_inp_bits_2(DecoupledStage_1_io_inp_bits_2),
    .io_inp_bits_3(DecoupledStage_1_io_inp_bits_3),
    .io_inp_bits_4(DecoupledStage_1_io_inp_bits_4),
    .io_inp_bits_5(DecoupledStage_1_io_inp_bits_5),
    .io_inp_bits_6(DecoupledStage_1_io_inp_bits_6),
    .io_inp_bits_7(DecoupledStage_1_io_inp_bits_7),
    .io_out_ready(DecoupledStage_1_io_out_ready),
    .io_out_valid(DecoupledStage_1_io_out_valid),
    .io_out_bits_0(DecoupledStage_1_io_out_bits_0),
    .io_out_bits_1(DecoupledStage_1_io_out_bits_1),
    .io_out_bits_2(DecoupledStage_1_io_out_bits_2),
    .io_out_bits_3(DecoupledStage_1_io_out_bits_3),
    .io_out_bits_4(DecoupledStage_1_io_out_bits_4),
    .io_out_bits_5(DecoupledStage_1_io_out_bits_5),
    .io_out_bits_6(DecoupledStage_1_io_out_bits_6),
    .io_out_bits_7(DecoupledStage_1_io_out_bits_7)
  );
  Queue_1 Queue ( // @[Decoupled.scala 294:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_0(Queue_io_enq_bits_0),
    .io_enq_bits_1(Queue_io_enq_bits_1),
    .io_enq_bits_2(Queue_io_enq_bits_2),
    .io_enq_bits_3(Queue_io_enq_bits_3),
    .io_enq_bits_4(Queue_io_enq_bits_4),
    .io_enq_bits_5(Queue_io_enq_bits_5),
    .io_enq_bits_6(Queue_io_enq_bits_6),
    .io_enq_bits_7(Queue_io_enq_bits_7),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_0(Queue_io_deq_bits_0),
    .io_deq_bits_1(Queue_io_deq_bits_1),
    .io_deq_bits_2(Queue_io_deq_bits_2),
    .io_deq_bits_3(Queue_io_deq_bits_3),
    .io_deq_bits_4(Queue_io_deq_bits_4),
    .io_deq_bits_5(Queue_io_deq_bits_5),
    .io_deq_bits_6(Queue_io_deq_bits_6),
    .io_deq_bits_7(Queue_io_deq_bits_7)
  );
  Queue_2 Queue_1 ( // @[Decoupled.scala 294:21]
    .clock(Queue_1_clock),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits_0(Queue_1_io_enq_bits_0),
    .io_enq_bits_1(Queue_1_io_enq_bits_1),
    .io_enq_bits_2(Queue_1_io_enq_bits_2),
    .io_enq_bits_3(Queue_1_io_enq_bits_3),
    .io_enq_bits_4(Queue_1_io_enq_bits_4),
    .io_enq_bits_5(Queue_1_io_enq_bits_5),
    .io_enq_bits_6(Queue_1_io_enq_bits_6),
    .io_enq_bits_7(Queue_1_io_enq_bits_7),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits_0(Queue_1_io_deq_bits_0),
    .io_deq_bits_1(Queue_1_io_deq_bits_1),
    .io_deq_bits_2(Queue_1_io_deq_bits_2),
    .io_deq_bits_3(Queue_1_io_deq_bits_3),
    .io_deq_bits_4(Queue_1_io_deq_bits_4),
    .io_deq_bits_5(Queue_1_io_deq_bits_5),
    .io_deq_bits_6(Queue_1_io_deq_bits_6),
    .io_deq_bits_7(Queue_1_io_deq_bits_7)
  );
  DecoupledStage DecoupledStage_2 ( // @[DecoupledStage.scala 30:19]
    .clock(DecoupledStage_2_clock),
    .reset(DecoupledStage_2_reset),
    .io_inp_ready(DecoupledStage_2_io_inp_ready),
    .io_inp_valid(DecoupledStage_2_io_inp_valid),
    .io_inp_bits_0(DecoupledStage_2_io_inp_bits_0),
    .io_inp_bits_1(DecoupledStage_2_io_inp_bits_1),
    .io_inp_bits_2(DecoupledStage_2_io_inp_bits_2),
    .io_inp_bits_3(DecoupledStage_2_io_inp_bits_3),
    .io_inp_bits_4(DecoupledStage_2_io_inp_bits_4),
    .io_inp_bits_5(DecoupledStage_2_io_inp_bits_5),
    .io_inp_bits_6(DecoupledStage_2_io_inp_bits_6),
    .io_inp_bits_7(DecoupledStage_2_io_inp_bits_7),
    .io_out_ready(DecoupledStage_2_io_out_ready),
    .io_out_valid(DecoupledStage_2_io_out_valid),
    .io_out_bits_0(DecoupledStage_2_io_out_bits_0),
    .io_out_bits_1(DecoupledStage_2_io_out_bits_1),
    .io_out_bits_2(DecoupledStage_2_io_out_bits_2),
    .io_out_bits_3(DecoupledStage_2_io_out_bits_3),
    .io_out_bits_4(DecoupledStage_2_io_out_bits_4),
    .io_out_bits_5(DecoupledStage_2_io_out_bits_5),
    .io_out_bits_6(DecoupledStage_2_io_out_bits_6),
    .io_out_bits_7(DecoupledStage_2_io_out_bits_7)
  );
  DecoupledStage DecoupledStage_3 ( // @[DecoupledStage.scala 30:19]
    .clock(DecoupledStage_3_clock),
    .reset(DecoupledStage_3_reset),
    .io_inp_ready(DecoupledStage_3_io_inp_ready),
    .io_inp_valid(DecoupledStage_3_io_inp_valid),
    .io_inp_bits_0(DecoupledStage_3_io_inp_bits_0),
    .io_inp_bits_1(DecoupledStage_3_io_inp_bits_1),
    .io_inp_bits_2(DecoupledStage_3_io_inp_bits_2),
    .io_inp_bits_3(DecoupledStage_3_io_inp_bits_3),
    .io_inp_bits_4(DecoupledStage_3_io_inp_bits_4),
    .io_inp_bits_5(DecoupledStage_3_io_inp_bits_5),
    .io_inp_bits_6(DecoupledStage_3_io_inp_bits_6),
    .io_inp_bits_7(DecoupledStage_3_io_inp_bits_7),
    .io_out_ready(DecoupledStage_3_io_out_ready),
    .io_out_valid(DecoupledStage_3_io_out_valid),
    .io_out_bits_0(DecoupledStage_3_io_out_bits_0),
    .io_out_bits_1(DecoupledStage_3_io_out_bits_1),
    .io_out_bits_2(DecoupledStage_3_io_out_bits_2),
    .io_out_bits_3(DecoupledStage_3_io_out_bits_3),
    .io_out_bits_4(DecoupledStage_3_io_out_bits_4),
    .io_out_bits_5(DecoupledStage_3_io_out_bits_5),
    .io_out_bits_6(DecoupledStage_3_io_out_bits_6),
    .io_out_bits_7(DecoupledStage_3_io_out_bits_7)
  );
  DecoupledStage_2 DecoupledStage_4 ( // @[DecoupledStage.scala 30:19]
    .clock(DecoupledStage_4_clock),
    .reset(DecoupledStage_4_reset),
    .io_inp_ready(DecoupledStage_4_io_inp_ready),
    .io_inp_valid(DecoupledStage_4_io_inp_valid),
    .io_inp_bits_0(DecoupledStage_4_io_inp_bits_0),
    .io_inp_bits_1(DecoupledStage_4_io_inp_bits_1),
    .io_inp_bits_2(DecoupledStage_4_io_inp_bits_2),
    .io_inp_bits_3(DecoupledStage_4_io_inp_bits_3),
    .io_inp_bits_4(DecoupledStage_4_io_inp_bits_4),
    .io_inp_bits_5(DecoupledStage_4_io_inp_bits_5),
    .io_inp_bits_6(DecoupledStage_4_io_inp_bits_6),
    .io_inp_bits_7(DecoupledStage_4_io_inp_bits_7),
    .io_out_ready(DecoupledStage_4_io_out_ready),
    .io_out_valid(DecoupledStage_4_io_out_valid),
    .io_out_bits_0(DecoupledStage_4_io_out_bits_0),
    .io_out_bits_1(DecoupledStage_4_io_out_bits_1),
    .io_out_bits_2(DecoupledStage_4_io_out_bits_2),
    .io_out_bits_3(DecoupledStage_4_io_out_bits_3),
    .io_out_bits_4(DecoupledStage_4_io_out_bits_4),
    .io_out_bits_5(DecoupledStage_4_io_out_bits_5),
    .io_out_bits_6(DecoupledStage_4_io_out_bits_6),
    .io_out_bits_7(DecoupledStage_4_io_out_bits_7)
  );
  assign _T = io_modeCompute == 1'h0; // @[trws.scala 68:16]
  assign _T_1 = _T | backend_io_done; // @[trws.scala 68:32]
  assign _T_2 = io_modeLoad == 1'h0; // @[trws.scala 68:57]
  assign _T_3 = _T_2 | loaf_io_doneLoading; // @[trws.scala 68:70]
  assign io_done = _T_1 & _T_3; // @[trws.scala 68:11]
  assign io_gi_ready = frontend_io_gi_ready; // @[trws.scala 46:18]
  assign io_wi_ready = frontend_io_wi_ready; // @[trws.scala 47:18]
  assign io_mi_ready = splitter_io_mi_ready; // @[trws.scala 38:18]
  assign io_slc_ready = loaf_io_slc_ready; // @[trws.scala 52:15]
  assign io_lof_ready = loaf_io_lof_ready; // @[trws.scala 53:15]
  assign io_mo_valid = backend_io_mo_valid; // @[trws.scala 67:9]
  assign io_mo_bits_bits_0 = backend_io_mo_bits_bits_0; // @[trws.scala 67:9]
  assign io_mo_bits_bits_1 = backend_io_mo_bits_bits_1; // @[trws.scala 67:9]
  assign io_mo_bits_bits_2 = backend_io_mo_bits_bits_2; // @[trws.scala 67:9]
  assign io_mo_bits_bits_3 = backend_io_mo_bits_bits_3; // @[trws.scala 67:9]
  assign io_mo_bits_bits_4 = backend_io_mo_bits_bits_4; // @[trws.scala 67:9]
  assign io_mo_bits_bits_5 = backend_io_mo_bits_bits_5; // @[trws.scala 67:9]
  assign io_mo_bits_bits_6 = backend_io_mo_bits_bits_6; // @[trws.scala 67:9]
  assign io_mo_bits_bits_7 = backend_io_mo_bits_bits_7; // @[trws.scala 67:9]
  assign splitter_io_mi_valid = io_mi_valid; // @[trws.scala 38:18]
  assign splitter_io_mi_bits_0 = io_mi_bits_0; // @[trws.scala 38:18]
  assign splitter_io_mi_bits_1 = io_mi_bits_1; // @[trws.scala 38:18]
  assign splitter_io_mi_bits_2 = io_mi_bits_2; // @[trws.scala 38:18]
  assign splitter_io_mi_bits_3 = io_mi_bits_3; // @[trws.scala 38:18]
  assign splitter_io_mi_bits_4 = io_mi_bits_4; // @[trws.scala 38:18]
  assign splitter_io_mi_bits_5 = io_mi_bits_5; // @[trws.scala 38:18]
  assign splitter_io_mi_bits_6 = io_mi_bits_6; // @[trws.scala 38:18]
  assign splitter_io_mi_bits_7 = io_mi_bits_7; // @[trws.scala 38:18]
  assign splitter_io_mi0_ready = DecoupledStage_io_inp_ready; // @[DecoupledStage.scala 33:15]
  assign splitter_io_mi1_ready = Queue_io_enq_ready; // @[Decoupled.scala 297:17]
  assign frontend_clock = clock;
  assign frontend_reset = reset;
  assign frontend_io_start = io_start; // @[trws.scala 49:21]
  assign frontend_io_gi_valid = io_gi_valid; // @[trws.scala 46:18]
  assign frontend_io_gi_bits_0 = io_gi_bits_0; // @[trws.scala 46:18]
  assign frontend_io_gi_bits_1 = io_gi_bits_1; // @[trws.scala 46:18]
  assign frontend_io_gi_bits_2 = io_gi_bits_2; // @[trws.scala 46:18]
  assign frontend_io_gi_bits_3 = io_gi_bits_3; // @[trws.scala 46:18]
  assign frontend_io_gi_bits_4 = io_gi_bits_4; // @[trws.scala 46:18]
  assign frontend_io_gi_bits_5 = io_gi_bits_5; // @[trws.scala 46:18]
  assign frontend_io_gi_bits_6 = io_gi_bits_6; // @[trws.scala 46:18]
  assign frontend_io_gi_bits_7 = io_gi_bits_7; // @[trws.scala 46:18]
  assign frontend_io_wi_valid = io_wi_valid; // @[trws.scala 47:18]
  assign frontend_io_wi_bits_0 = io_wi_bits_0; // @[trws.scala 47:18]
  assign frontend_io_wi_bits_1 = io_wi_bits_1; // @[trws.scala 47:18]
  assign frontend_io_wi_bits_2 = io_wi_bits_2; // @[trws.scala 47:18]
  assign frontend_io_wi_bits_3 = io_wi_bits_3; // @[trws.scala 47:18]
  assign frontend_io_wi_bits_4 = io_wi_bits_4; // @[trws.scala 47:18]
  assign frontend_io_wi_bits_5 = io_wi_bits_5; // @[trws.scala 47:18]
  assign frontend_io_wi_bits_6 = io_wi_bits_6; // @[trws.scala 47:18]
  assign frontend_io_wi_bits_7 = io_wi_bits_7; // @[trws.scala 47:18]
  assign frontend_io_a0_valid = DecoupledStage_1_io_out_valid; // @[trws.scala 44:18]
  assign frontend_io_a0_bits_0 = DecoupledStage_1_io_out_bits_0; // @[trws.scala 44:18]
  assign frontend_io_a0_bits_1 = DecoupledStage_1_io_out_bits_1; // @[trws.scala 44:18]
  assign frontend_io_a0_bits_2 = DecoupledStage_1_io_out_bits_2; // @[trws.scala 44:18]
  assign frontend_io_a0_bits_3 = DecoupledStage_1_io_out_bits_3; // @[trws.scala 44:18]
  assign frontend_io_a0_bits_4 = DecoupledStage_1_io_out_bits_4; // @[trws.scala 44:18]
  assign frontend_io_a0_bits_5 = DecoupledStage_1_io_out_bits_5; // @[trws.scala 44:18]
  assign frontend_io_a0_bits_6 = DecoupledStage_1_io_out_bits_6; // @[trws.scala 44:18]
  assign frontend_io_a0_bits_7 = DecoupledStage_1_io_out_bits_7; // @[trws.scala 44:18]
  assign frontend_io_mi1_valid = Queue_io_deq_valid; // @[trws.scala 45:19]
  assign frontend_io_mi1_bits_0 = Queue_io_deq_bits_0; // @[trws.scala 45:19]
  assign frontend_io_mi1_bits_1 = Queue_io_deq_bits_1; // @[trws.scala 45:19]
  assign frontend_io_mi1_bits_2 = Queue_io_deq_bits_2; // @[trws.scala 45:19]
  assign frontend_io_mi1_bits_3 = Queue_io_deq_bits_3; // @[trws.scala 45:19]
  assign frontend_io_mi1_bits_4 = Queue_io_deq_bits_4; // @[trws.scala 45:19]
  assign frontend_io_mi1_bits_5 = Queue_io_deq_bits_5; // @[trws.scala 45:19]
  assign frontend_io_mi1_bits_6 = Queue_io_deq_bits_6; // @[trws.scala 45:19]
  assign frontend_io_mi1_bits_7 = Queue_io_deq_bits_7; // @[trws.scala 45:19]
  assign frontend_io_adj_valid = Queue_1_io_deq_valid; // @[trws.scala 48:19]
  assign frontend_io_adj_bits_0 = Queue_1_io_deq_bits_0; // @[trws.scala 48:19]
  assign frontend_io_adj_bits_1 = Queue_1_io_deq_bits_1; // @[trws.scala 48:19]
  assign frontend_io_adj_bits_2 = Queue_1_io_deq_bits_2; // @[trws.scala 48:19]
  assign frontend_io_adj_bits_3 = Queue_1_io_deq_bits_3; // @[trws.scala 48:19]
  assign frontend_io_adj_bits_4 = Queue_1_io_deq_bits_4; // @[trws.scala 48:19]
  assign frontend_io_adj_bits_5 = Queue_1_io_deq_bits_5; // @[trws.scala 48:19]
  assign frontend_io_adj_bits_6 = Queue_1_io_deq_bits_6; // @[trws.scala 48:19]
  assign frontend_io_adj_bits_7 = Queue_1_io_deq_bits_7; // @[trws.scala 48:19]
  assign frontend_io_off_ready = DecoupledStage_2_io_inp_ready; // @[DecoupledStage.scala 33:15]
  assign backend_clock = clock;
  assign backend_reset = reset;
  assign backend_io_start = io_start; // @[trws.scala 65:20]
  assign backend_io_res_valid = DecoupledStage_4_io_out_valid; // @[trws.scala 64:18]
  assign backend_io_res_bits_0 = DecoupledStage_4_io_out_bits_0; // @[trws.scala 64:18]
  assign backend_io_res_bits_1 = DecoupledStage_4_io_out_bits_1; // @[trws.scala 64:18]
  assign backend_io_res_bits_2 = DecoupledStage_4_io_out_bits_2; // @[trws.scala 64:18]
  assign backend_io_res_bits_3 = DecoupledStage_4_io_out_bits_3; // @[trws.scala 64:18]
  assign backend_io_res_bits_4 = DecoupledStage_4_io_out_bits_4; // @[trws.scala 64:18]
  assign backend_io_res_bits_5 = DecoupledStage_4_io_out_bits_5; // @[trws.scala 64:18]
  assign backend_io_res_bits_6 = DecoupledStage_4_io_out_bits_6; // @[trws.scala 64:18]
  assign backend_io_res_bits_7 = DecoupledStage_4_io_out_bits_7; // @[trws.scala 64:18]
  assign backend_io_mo_ready = io_mo_ready; // @[trws.scala 67:9]
  assign backend_io_adj_ready = Queue_1_io_enq_ready; // @[Decoupled.scala 297:17]
  assign accumulator_clock = clock;
  assign accumulator_reset = reset;
  assign accumulator_io_mi0_valid = DecoupledStage_io_out_valid; // @[trws.scala 41:22]
  assign accumulator_io_mi0_bits_0 = DecoupledStage_io_out_bits_0; // @[trws.scala 41:22]
  assign accumulator_io_mi0_bits_1 = DecoupledStage_io_out_bits_1; // @[trws.scala 41:22]
  assign accumulator_io_mi0_bits_2 = DecoupledStage_io_out_bits_2; // @[trws.scala 41:22]
  assign accumulator_io_mi0_bits_3 = DecoupledStage_io_out_bits_3; // @[trws.scala 41:22]
  assign accumulator_io_mi0_bits_4 = DecoupledStage_io_out_bits_4; // @[trws.scala 41:22]
  assign accumulator_io_mi0_bits_5 = DecoupledStage_io_out_bits_5; // @[trws.scala 41:22]
  assign accumulator_io_mi0_bits_6 = DecoupledStage_io_out_bits_6; // @[trws.scala 41:22]
  assign accumulator_io_mi0_bits_7 = DecoupledStage_io_out_bits_7; // @[trws.scala 41:22]
  assign accumulator_io_a0_ready = DecoupledStage_1_io_inp_ready; // @[DecoupledStage.scala 33:15]
  assign loaf_clock = clock;
  assign loaf_reset = reset;
  assign loaf_io_start = io_start; // @[trws.scala 55:17]
  assign loaf_io_modeLoad = io_modeLoad; // @[trws.scala 56:20]
  assign loaf_io_modeCompute = io_modeCompute; // @[trws.scala 57:23]
  assign loaf_io_loadIdx = io_loadIdx; // @[trws.scala 58:19]
  assign loaf_io_computeIdx = io_computeIdx; // @[trws.scala 59:22]
  assign loaf_io_off_valid = DecoupledStage_2_io_out_valid; // @[trws.scala 51:15]
  assign loaf_io_off_bits_0 = DecoupledStage_2_io_out_bits_0; // @[trws.scala 51:15]
  assign loaf_io_off_bits_1 = DecoupledStage_2_io_out_bits_1; // @[trws.scala 51:15]
  assign loaf_io_off_bits_2 = DecoupledStage_2_io_out_bits_2; // @[trws.scala 51:15]
  assign loaf_io_off_bits_3 = DecoupledStage_2_io_out_bits_3; // @[trws.scala 51:15]
  assign loaf_io_off_bits_4 = DecoupledStage_2_io_out_bits_4; // @[trws.scala 51:15]
  assign loaf_io_off_bits_5 = DecoupledStage_2_io_out_bits_5; // @[trws.scala 51:15]
  assign loaf_io_off_bits_6 = DecoupledStage_2_io_out_bits_6; // @[trws.scala 51:15]
  assign loaf_io_off_bits_7 = DecoupledStage_2_io_out_bits_7; // @[trws.scala 51:15]
  assign loaf_io_out_ready = DecoupledStage_3_io_inp_ready; // @[DecoupledStage.scala 33:15]
  assign loaf_io_slc_valid = io_slc_valid; // @[trws.scala 52:15]
  assign loaf_io_slc_bits_e = io_slc_bits_e; // @[trws.scala 52:15]
  assign loaf_io_slc_bits_a = io_slc_bits_a; // @[trws.scala 52:15]
  assign loaf_io_lof_valid = io_lof_valid; // @[trws.scala 53:15]
  assign loaf_io_lof_bits_e = io_lof_bits_e; // @[trws.scala 53:15]
  assign loaf_io_lof_bits_a = io_lof_bits_a; // @[trws.scala 53:15]
  assign clamper_clock = clock;
  assign clamper_reset = reset;
  assign clamper_io_start = io_start; // @[trws.scala 62:20]
  assign clamper_io_out_valid = DecoupledStage_3_io_out_valid; // @[trws.scala 61:18]
  assign clamper_io_out_bits_0 = DecoupledStage_3_io_out_bits_0; // @[trws.scala 61:18]
  assign clamper_io_out_bits_1 = DecoupledStage_3_io_out_bits_1; // @[trws.scala 61:18]
  assign clamper_io_out_bits_2 = DecoupledStage_3_io_out_bits_2; // @[trws.scala 61:18]
  assign clamper_io_out_bits_3 = DecoupledStage_3_io_out_bits_3; // @[trws.scala 61:18]
  assign clamper_io_out_bits_4 = DecoupledStage_3_io_out_bits_4; // @[trws.scala 61:18]
  assign clamper_io_out_bits_5 = DecoupledStage_3_io_out_bits_5; // @[trws.scala 61:18]
  assign clamper_io_out_bits_6 = DecoupledStage_3_io_out_bits_6; // @[trws.scala 61:18]
  assign clamper_io_out_bits_7 = DecoupledStage_3_io_out_bits_7; // @[trws.scala 61:18]
  assign clamper_io_res_ready = DecoupledStage_4_io_inp_ready; // @[DecoupledStage.scala 33:15]
  assign DecoupledStage_clock = clock;
  assign DecoupledStage_reset = reset;
  assign DecoupledStage_io_inp_valid = splitter_io_mi0_valid; // @[DecoupledStage.scala 31:20]
  assign DecoupledStage_io_inp_bits_0 = splitter_io_mi0_bits_0; // @[DecoupledStage.scala 32:19]
  assign DecoupledStage_io_inp_bits_1 = splitter_io_mi0_bits_1; // @[DecoupledStage.scala 32:19]
  assign DecoupledStage_io_inp_bits_2 = splitter_io_mi0_bits_2; // @[DecoupledStage.scala 32:19]
  assign DecoupledStage_io_inp_bits_3 = splitter_io_mi0_bits_3; // @[DecoupledStage.scala 32:19]
  assign DecoupledStage_io_inp_bits_4 = splitter_io_mi0_bits_4; // @[DecoupledStage.scala 32:19]
  assign DecoupledStage_io_inp_bits_5 = splitter_io_mi0_bits_5; // @[DecoupledStage.scala 32:19]
  assign DecoupledStage_io_inp_bits_6 = splitter_io_mi0_bits_6; // @[DecoupledStage.scala 32:19]
  assign DecoupledStage_io_inp_bits_7 = splitter_io_mi0_bits_7; // @[DecoupledStage.scala 32:19]
  assign DecoupledStage_io_out_ready = accumulator_io_mi0_ready; // @[trws.scala 41:22]
  assign DecoupledStage_1_clock = clock;
  assign DecoupledStage_1_reset = reset;
  assign DecoupledStage_1_io_inp_valid = accumulator_io_a0_valid; // @[DecoupledStage.scala 31:20]
  assign DecoupledStage_1_io_inp_bits_0 = accumulator_io_a0_bits_0; // @[DecoupledStage.scala 32:19]
  assign DecoupledStage_1_io_inp_bits_1 = accumulator_io_a0_bits_1; // @[DecoupledStage.scala 32:19]
  assign DecoupledStage_1_io_inp_bits_2 = accumulator_io_a0_bits_2; // @[DecoupledStage.scala 32:19]
  assign DecoupledStage_1_io_inp_bits_3 = accumulator_io_a0_bits_3; // @[DecoupledStage.scala 32:19]
  assign DecoupledStage_1_io_inp_bits_4 = accumulator_io_a0_bits_4; // @[DecoupledStage.scala 32:19]
  assign DecoupledStage_1_io_inp_bits_5 = accumulator_io_a0_bits_5; // @[DecoupledStage.scala 32:19]
  assign DecoupledStage_1_io_inp_bits_6 = accumulator_io_a0_bits_6; // @[DecoupledStage.scala 32:19]
  assign DecoupledStage_1_io_inp_bits_7 = accumulator_io_a0_bits_7; // @[DecoupledStage.scala 32:19]
  assign DecoupledStage_1_io_out_ready = frontend_io_a0_ready; // @[trws.scala 44:18]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = splitter_io_mi1_valid; // @[Decoupled.scala 295:22]
  assign Queue_io_enq_bits_0 = splitter_io_mi1_bits_0; // @[Decoupled.scala 296:21]
  assign Queue_io_enq_bits_1 = splitter_io_mi1_bits_1; // @[Decoupled.scala 296:21]
  assign Queue_io_enq_bits_2 = splitter_io_mi1_bits_2; // @[Decoupled.scala 296:21]
  assign Queue_io_enq_bits_3 = splitter_io_mi1_bits_3; // @[Decoupled.scala 296:21]
  assign Queue_io_enq_bits_4 = splitter_io_mi1_bits_4; // @[Decoupled.scala 296:21]
  assign Queue_io_enq_bits_5 = splitter_io_mi1_bits_5; // @[Decoupled.scala 296:21]
  assign Queue_io_enq_bits_6 = splitter_io_mi1_bits_6; // @[Decoupled.scala 296:21]
  assign Queue_io_enq_bits_7 = splitter_io_mi1_bits_7; // @[Decoupled.scala 296:21]
  assign Queue_io_deq_ready = frontend_io_mi1_ready; // @[trws.scala 45:19]
  assign Queue_1_clock = clock;
  assign Queue_1_reset = reset;
  assign Queue_1_io_enq_valid = backend_io_adj_valid; // @[Decoupled.scala 295:22]
  assign Queue_1_io_enq_bits_0 = backend_io_adj_bits_0; // @[Decoupled.scala 296:21]
  assign Queue_1_io_enq_bits_1 = backend_io_adj_bits_1; // @[Decoupled.scala 296:21]
  assign Queue_1_io_enq_bits_2 = backend_io_adj_bits_2; // @[Decoupled.scala 296:21]
  assign Queue_1_io_enq_bits_3 = backend_io_adj_bits_3; // @[Decoupled.scala 296:21]
  assign Queue_1_io_enq_bits_4 = backend_io_adj_bits_4; // @[Decoupled.scala 296:21]
  assign Queue_1_io_enq_bits_5 = backend_io_adj_bits_5; // @[Decoupled.scala 296:21]
  assign Queue_1_io_enq_bits_6 = backend_io_adj_bits_6; // @[Decoupled.scala 296:21]
  assign Queue_1_io_enq_bits_7 = backend_io_adj_bits_7; // @[Decoupled.scala 296:21]
  assign Queue_1_io_deq_ready = frontend_io_adj_ready; // @[trws.scala 48:19]
  assign DecoupledStage_2_clock = clock;
  assign DecoupledStage_2_reset = reset;
  assign DecoupledStage_2_io_inp_valid = frontend_io_off_valid; // @[DecoupledStage.scala 31:20]
  assign DecoupledStage_2_io_inp_bits_0 = frontend_io_off_bits_0; // @[DecoupledStage.scala 32:19]
  assign DecoupledStage_2_io_inp_bits_1 = frontend_io_off_bits_1; // @[DecoupledStage.scala 32:19]
  assign DecoupledStage_2_io_inp_bits_2 = frontend_io_off_bits_2; // @[DecoupledStage.scala 32:19]
  assign DecoupledStage_2_io_inp_bits_3 = frontend_io_off_bits_3; // @[DecoupledStage.scala 32:19]
  assign DecoupledStage_2_io_inp_bits_4 = frontend_io_off_bits_4; // @[DecoupledStage.scala 32:19]
  assign DecoupledStage_2_io_inp_bits_5 = frontend_io_off_bits_5; // @[DecoupledStage.scala 32:19]
  assign DecoupledStage_2_io_inp_bits_6 = frontend_io_off_bits_6; // @[DecoupledStage.scala 32:19]
  assign DecoupledStage_2_io_inp_bits_7 = frontend_io_off_bits_7; // @[DecoupledStage.scala 32:19]
  assign DecoupledStage_2_io_out_ready = loaf_io_off_ready; // @[trws.scala 51:15]
  assign DecoupledStage_3_clock = clock;
  assign DecoupledStage_3_reset = reset;
  assign DecoupledStage_3_io_inp_valid = loaf_io_out_valid; // @[DecoupledStage.scala 31:20]
  assign DecoupledStage_3_io_inp_bits_0 = loaf_io_out_bits_0; // @[DecoupledStage.scala 32:19]
  assign DecoupledStage_3_io_inp_bits_1 = loaf_io_out_bits_1; // @[DecoupledStage.scala 32:19]
  assign DecoupledStage_3_io_inp_bits_2 = loaf_io_out_bits_2; // @[DecoupledStage.scala 32:19]
  assign DecoupledStage_3_io_inp_bits_3 = loaf_io_out_bits_3; // @[DecoupledStage.scala 32:19]
  assign DecoupledStage_3_io_inp_bits_4 = loaf_io_out_bits_4; // @[DecoupledStage.scala 32:19]
  assign DecoupledStage_3_io_inp_bits_5 = loaf_io_out_bits_5; // @[DecoupledStage.scala 32:19]
  assign DecoupledStage_3_io_inp_bits_6 = loaf_io_out_bits_6; // @[DecoupledStage.scala 32:19]
  assign DecoupledStage_3_io_inp_bits_7 = loaf_io_out_bits_7; // @[DecoupledStage.scala 32:19]
  assign DecoupledStage_3_io_out_ready = clamper_io_out_ready; // @[trws.scala 61:18]
  assign DecoupledStage_4_clock = clock;
  assign DecoupledStage_4_reset = reset;
  assign DecoupledStage_4_io_inp_valid = clamper_io_res_valid; // @[DecoupledStage.scala 31:20]
  assign DecoupledStage_4_io_inp_bits_0 = clamper_io_res_bits_0; // @[DecoupledStage.scala 32:19]
  assign DecoupledStage_4_io_inp_bits_1 = clamper_io_res_bits_1; // @[DecoupledStage.scala 32:19]
  assign DecoupledStage_4_io_inp_bits_2 = clamper_io_res_bits_2; // @[DecoupledStage.scala 32:19]
  assign DecoupledStage_4_io_inp_bits_3 = clamper_io_res_bits_3; // @[DecoupledStage.scala 32:19]
  assign DecoupledStage_4_io_inp_bits_4 = clamper_io_res_bits_4; // @[DecoupledStage.scala 32:19]
  assign DecoupledStage_4_io_inp_bits_5 = clamper_io_res_bits_5; // @[DecoupledStage.scala 32:19]
  assign DecoupledStage_4_io_inp_bits_6 = clamper_io_res_bits_6; // @[DecoupledStage.scala 32:19]
  assign DecoupledStage_4_io_inp_bits_7 = clamper_io_res_bits_7; // @[DecoupledStage.scala 32:19]
  assign DecoupledStage_4_io_out_ready = backend_io_res_ready; // @[trws.scala 64:18]
endmodule
module trwsWrapper(
  input         clock,
  input         reset,
  input         io_start,
  output        io_done,
  input         io_modeLoad,
  input         io_modeCompute,
  input         io_loadIdx,
  input         io_computeIdx,
  output        io_gi_ready,
  input         io_gi_valid,
  input  [15:0] io_gi_bits_0,
  input  [15:0] io_gi_bits_1,
  input  [15:0] io_gi_bits_2,
  input  [15:0] io_gi_bits_3,
  input  [15:0] io_gi_bits_4,
  input  [15:0] io_gi_bits_5,
  input  [15:0] io_gi_bits_6,
  input  [15:0] io_gi_bits_7,
  output        io_wi_ready,
  input         io_wi_valid,
  input  [15:0] io_wi_bits_0,
  input  [15:0] io_wi_bits_1,
  input  [15:0] io_wi_bits_2,
  input  [15:0] io_wi_bits_3,
  input  [15:0] io_wi_bits_4,
  input  [15:0] io_wi_bits_5,
  input  [15:0] io_wi_bits_6,
  input  [15:0] io_wi_bits_7,
  output        io_mi_ready,
  input         io_mi_valid,
  input  [15:0] io_mi_bits_0,
  input  [15:0] io_mi_bits_1,
  input  [15:0] io_mi_bits_2,
  input  [15:0] io_mi_bits_3,
  input  [15:0] io_mi_bits_4,
  input  [15:0] io_mi_bits_5,
  input  [15:0] io_mi_bits_6,
  input  [15:0] io_mi_bits_7,
  output        io_slc_ready,
  input         io_slc_valid,
  input  [15:0] io_slc_bits_e,
  input  [15:0] io_slc_bits_a,
  output        io_lof_ready,
  input         io_lof_valid,
  input  [15:0] io_lof_bits_e,
  input  [15:0] io_lof_bits_a,
  input         io_mo_ready,
  output        io_mo_valid,
  output [15:0] io_mo_bits_0,
  output [15:0] io_mo_bits_1,
  output [15:0] io_mo_bits_2,
  output [15:0] io_mo_bits_3,
  output [15:0] io_mo_bits_4,
  output [15:0] io_mo_bits_5,
  output [15:0] io_mo_bits_6,
  output [15:0] io_mo_bits_7
);
  wire  m_clock; // @[trws.scala 93:17]
  wire  m_reset; // @[trws.scala 93:17]
  wire  m_io_start; // @[trws.scala 93:17]
  wire  m_io_done; // @[trws.scala 93:17]
  wire  m_io_modeLoad; // @[trws.scala 93:17]
  wire  m_io_modeCompute; // @[trws.scala 93:17]
  wire  m_io_loadIdx; // @[trws.scala 93:17]
  wire  m_io_computeIdx; // @[trws.scala 93:17]
  wire  m_io_gi_ready; // @[trws.scala 93:17]
  wire  m_io_gi_valid; // @[trws.scala 93:17]
  wire [15:0] m_io_gi_bits_0; // @[trws.scala 93:17]
  wire [15:0] m_io_gi_bits_1; // @[trws.scala 93:17]
  wire [15:0] m_io_gi_bits_2; // @[trws.scala 93:17]
  wire [15:0] m_io_gi_bits_3; // @[trws.scala 93:17]
  wire [15:0] m_io_gi_bits_4; // @[trws.scala 93:17]
  wire [15:0] m_io_gi_bits_5; // @[trws.scala 93:17]
  wire [15:0] m_io_gi_bits_6; // @[trws.scala 93:17]
  wire [15:0] m_io_gi_bits_7; // @[trws.scala 93:17]
  wire  m_io_wi_ready; // @[trws.scala 93:17]
  wire  m_io_wi_valid; // @[trws.scala 93:17]
  wire [15:0] m_io_wi_bits_0; // @[trws.scala 93:17]
  wire [15:0] m_io_wi_bits_1; // @[trws.scala 93:17]
  wire [15:0] m_io_wi_bits_2; // @[trws.scala 93:17]
  wire [15:0] m_io_wi_bits_3; // @[trws.scala 93:17]
  wire [15:0] m_io_wi_bits_4; // @[trws.scala 93:17]
  wire [15:0] m_io_wi_bits_5; // @[trws.scala 93:17]
  wire [15:0] m_io_wi_bits_6; // @[trws.scala 93:17]
  wire [15:0] m_io_wi_bits_7; // @[trws.scala 93:17]
  wire  m_io_mi_ready; // @[trws.scala 93:17]
  wire  m_io_mi_valid; // @[trws.scala 93:17]
  wire [15:0] m_io_mi_bits_0; // @[trws.scala 93:17]
  wire [15:0] m_io_mi_bits_1; // @[trws.scala 93:17]
  wire [15:0] m_io_mi_bits_2; // @[trws.scala 93:17]
  wire [15:0] m_io_mi_bits_3; // @[trws.scala 93:17]
  wire [15:0] m_io_mi_bits_4; // @[trws.scala 93:17]
  wire [15:0] m_io_mi_bits_5; // @[trws.scala 93:17]
  wire [15:0] m_io_mi_bits_6; // @[trws.scala 93:17]
  wire [15:0] m_io_mi_bits_7; // @[trws.scala 93:17]
  wire  m_io_slc_ready; // @[trws.scala 93:17]
  wire  m_io_slc_valid; // @[trws.scala 93:17]
  wire [15:0] m_io_slc_bits_e; // @[trws.scala 93:17]
  wire [15:0] m_io_slc_bits_a; // @[trws.scala 93:17]
  wire  m_io_lof_ready; // @[trws.scala 93:17]
  wire  m_io_lof_valid; // @[trws.scala 93:17]
  wire [15:0] m_io_lof_bits_e; // @[trws.scala 93:17]
  wire [15:0] m_io_lof_bits_a; // @[trws.scala 93:17]
  wire  m_io_mo_ready; // @[trws.scala 93:17]
  wire  m_io_mo_valid; // @[trws.scala 93:17]
  wire [15:0] m_io_mo_bits_bits_0; // @[trws.scala 93:17]
  wire [15:0] m_io_mo_bits_bits_1; // @[trws.scala 93:17]
  wire [15:0] m_io_mo_bits_bits_2; // @[trws.scala 93:17]
  wire [15:0] m_io_mo_bits_bits_3; // @[trws.scala 93:17]
  wire [15:0] m_io_mo_bits_bits_4; // @[trws.scala 93:17]
  wire [15:0] m_io_mo_bits_bits_5; // @[trws.scala 93:17]
  wire [15:0] m_io_mo_bits_bits_6; // @[trws.scala 93:17]
  wire [15:0] m_io_mo_bits_bits_7; // @[trws.scala 93:17]
  trws m ( // @[trws.scala 93:17]
    .clock(m_clock),
    .reset(m_reset),
    .io_start(m_io_start),
    .io_done(m_io_done),
    .io_modeLoad(m_io_modeLoad),
    .io_modeCompute(m_io_modeCompute),
    .io_loadIdx(m_io_loadIdx),
    .io_computeIdx(m_io_computeIdx),
    .io_gi_ready(m_io_gi_ready),
    .io_gi_valid(m_io_gi_valid),
    .io_gi_bits_0(m_io_gi_bits_0),
    .io_gi_bits_1(m_io_gi_bits_1),
    .io_gi_bits_2(m_io_gi_bits_2),
    .io_gi_bits_3(m_io_gi_bits_3),
    .io_gi_bits_4(m_io_gi_bits_4),
    .io_gi_bits_5(m_io_gi_bits_5),
    .io_gi_bits_6(m_io_gi_bits_6),
    .io_gi_bits_7(m_io_gi_bits_7),
    .io_wi_ready(m_io_wi_ready),
    .io_wi_valid(m_io_wi_valid),
    .io_wi_bits_0(m_io_wi_bits_0),
    .io_wi_bits_1(m_io_wi_bits_1),
    .io_wi_bits_2(m_io_wi_bits_2),
    .io_wi_bits_3(m_io_wi_bits_3),
    .io_wi_bits_4(m_io_wi_bits_4),
    .io_wi_bits_5(m_io_wi_bits_5),
    .io_wi_bits_6(m_io_wi_bits_6),
    .io_wi_bits_7(m_io_wi_bits_7),
    .io_mi_ready(m_io_mi_ready),
    .io_mi_valid(m_io_mi_valid),
    .io_mi_bits_0(m_io_mi_bits_0),
    .io_mi_bits_1(m_io_mi_bits_1),
    .io_mi_bits_2(m_io_mi_bits_2),
    .io_mi_bits_3(m_io_mi_bits_3),
    .io_mi_bits_4(m_io_mi_bits_4),
    .io_mi_bits_5(m_io_mi_bits_5),
    .io_mi_bits_6(m_io_mi_bits_6),
    .io_mi_bits_7(m_io_mi_bits_7),
    .io_slc_ready(m_io_slc_ready),
    .io_slc_valid(m_io_slc_valid),
    .io_slc_bits_e(m_io_slc_bits_e),
    .io_slc_bits_a(m_io_slc_bits_a),
    .io_lof_ready(m_io_lof_ready),
    .io_lof_valid(m_io_lof_valid),
    .io_lof_bits_e(m_io_lof_bits_e),
    .io_lof_bits_a(m_io_lof_bits_a),
    .io_mo_ready(m_io_mo_ready),
    .io_mo_valid(m_io_mo_valid),
    .io_mo_bits_bits_0(m_io_mo_bits_bits_0),
    .io_mo_bits_bits_1(m_io_mo_bits_bits_1),
    .io_mo_bits_bits_2(m_io_mo_bits_bits_2),
    .io_mo_bits_bits_3(m_io_mo_bits_bits_3),
    .io_mo_bits_bits_4(m_io_mo_bits_bits_4),
    .io_mo_bits_bits_5(m_io_mo_bits_bits_5),
    .io_mo_bits_bits_6(m_io_mo_bits_bits_6),
    .io_mo_bits_bits_7(m_io_mo_bits_bits_7)
  );
  assign io_done = m_io_done; // @[trws.scala 95:11]
  assign io_gi_ready = m_io_gi_ready; // @[trws.scala 103:11]
  assign io_wi_ready = m_io_wi_ready; // @[trws.scala 104:11]
  assign io_mi_ready = m_io_mi_ready; // @[trws.scala 105:11]
  assign io_slc_ready = m_io_slc_ready; // @[trws.scala 107:12]
  assign io_lof_ready = m_io_lof_ready; // @[trws.scala 108:12]
  assign io_mo_valid = m_io_mo_valid; // @[trws.scala 110:15]
  assign io_mo_bits_0 = m_io_mo_bits_bits_0; // @[trws.scala 111:14]
  assign io_mo_bits_1 = m_io_mo_bits_bits_1; // @[trws.scala 111:14]
  assign io_mo_bits_2 = m_io_mo_bits_bits_2; // @[trws.scala 111:14]
  assign io_mo_bits_3 = m_io_mo_bits_bits_3; // @[trws.scala 111:14]
  assign io_mo_bits_4 = m_io_mo_bits_bits_4; // @[trws.scala 111:14]
  assign io_mo_bits_5 = m_io_mo_bits_bits_5; // @[trws.scala 111:14]
  assign io_mo_bits_6 = m_io_mo_bits_bits_6; // @[trws.scala 111:14]
  assign io_mo_bits_7 = m_io_mo_bits_bits_7; // @[trws.scala 111:14]
  assign m_clock = clock;
  assign m_reset = reset;
  assign m_io_start = io_start; // @[trws.scala 94:14]
  assign m_io_modeLoad = io_modeLoad; // @[trws.scala 97:17]
  assign m_io_modeCompute = io_modeCompute; // @[trws.scala 98:20]
  assign m_io_loadIdx = io_loadIdx; // @[trws.scala 100:16]
  assign m_io_computeIdx = io_computeIdx; // @[trws.scala 101:19]
  assign m_io_gi_valid = io_gi_valid; // @[trws.scala 103:11]
  assign m_io_gi_bits_0 = io_gi_bits_0; // @[trws.scala 103:11]
  assign m_io_gi_bits_1 = io_gi_bits_1; // @[trws.scala 103:11]
  assign m_io_gi_bits_2 = io_gi_bits_2; // @[trws.scala 103:11]
  assign m_io_gi_bits_3 = io_gi_bits_3; // @[trws.scala 103:11]
  assign m_io_gi_bits_4 = io_gi_bits_4; // @[trws.scala 103:11]
  assign m_io_gi_bits_5 = io_gi_bits_5; // @[trws.scala 103:11]
  assign m_io_gi_bits_6 = io_gi_bits_6; // @[trws.scala 103:11]
  assign m_io_gi_bits_7 = io_gi_bits_7; // @[trws.scala 103:11]
  assign m_io_wi_valid = io_wi_valid; // @[trws.scala 104:11]
  assign m_io_wi_bits_0 = io_wi_bits_0; // @[trws.scala 104:11]
  assign m_io_wi_bits_1 = io_wi_bits_1; // @[trws.scala 104:11]
  assign m_io_wi_bits_2 = io_wi_bits_2; // @[trws.scala 104:11]
  assign m_io_wi_bits_3 = io_wi_bits_3; // @[trws.scala 104:11]
  assign m_io_wi_bits_4 = io_wi_bits_4; // @[trws.scala 104:11]
  assign m_io_wi_bits_5 = io_wi_bits_5; // @[trws.scala 104:11]
  assign m_io_wi_bits_6 = io_wi_bits_6; // @[trws.scala 104:11]
  assign m_io_wi_bits_7 = io_wi_bits_7; // @[trws.scala 104:11]
  assign m_io_mi_valid = io_mi_valid; // @[trws.scala 105:11]
  assign m_io_mi_bits_0 = io_mi_bits_0; // @[trws.scala 105:11]
  assign m_io_mi_bits_1 = io_mi_bits_1; // @[trws.scala 105:11]
  assign m_io_mi_bits_2 = io_mi_bits_2; // @[trws.scala 105:11]
  assign m_io_mi_bits_3 = io_mi_bits_3; // @[trws.scala 105:11]
  assign m_io_mi_bits_4 = io_mi_bits_4; // @[trws.scala 105:11]
  assign m_io_mi_bits_5 = io_mi_bits_5; // @[trws.scala 105:11]
  assign m_io_mi_bits_6 = io_mi_bits_6; // @[trws.scala 105:11]
  assign m_io_mi_bits_7 = io_mi_bits_7; // @[trws.scala 105:11]
  assign m_io_slc_valid = io_slc_valid; // @[trws.scala 107:12]
  assign m_io_slc_bits_e = io_slc_bits_e; // @[trws.scala 107:12]
  assign m_io_slc_bits_a = io_slc_bits_a; // @[trws.scala 107:12]
  assign m_io_lof_valid = io_lof_valid; // @[trws.scala 108:12]
  assign m_io_lof_bits_e = io_lof_bits_e; // @[trws.scala 108:12]
  assign m_io_lof_bits_a = io_lof_bits_a; // @[trws.scala 108:12]
  assign m_io_mo_ready = io_mo_ready; // @[trws.scala 113:17]
endmodule
